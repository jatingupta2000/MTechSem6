`timescale 1ns/10ps//time-unit = 1 ns and precision = 10 ps

module testbench ( );
  // Inputs
	reg v_in2_v;
  reg v_in3_v;
  reg v_in4_v;
  reg v_in5_v;
  reg v_in6_v;
  reg v_in7_v;
  reg v_in8_v;
  reg v_in9_v;
  reg v_in10_v;
  reg v_in11_v;
  reg v_in12_v;
  reg v_in13_v;
  reg v_in14_v;
  reg v_in15_v;
  reg v_in16_v;
  reg v_in17_v;
  reg v_in18_v;
  reg v_in19_v;
  reg v_in20_v;
  reg v_in21_v;
  reg v_in22_v;
  reg v_in23_v;
  reg v_in24_v;
  reg v_in25_v;
  reg v_in26_v;
  reg v_in27_v;
  reg v_in28_v;
  reg v_in29_v;
  reg v_in30_v;
  reg v_in31_v;
  reg v_in32_v;
  reg v_in33_v;
	reg v_keyinput_0_v;
	reg v_keyinput_1_v;
	reg v_keyinput_2_v;
	reg v_keyinput_3_v;
	reg v_keyinput_4_v;
	reg v_keyinput_5_v;
	reg v_keyinput_6_v;
	reg v_keyinput_7_v;
	reg v_keyinput_8_v;
	reg v_keyinput_9_v;
	reg v_keyinput_10_v;
	reg v_keyinput_11_v;
	reg v_keyinput_12_v;
	reg v_keyinput_13_v;
	reg v_keyinput_14_v;
	reg v_keyinput_15_v;
	reg v_keyinput_16_v;
	reg v_keyinput_17_v;
	reg v_keyinput_18_v;
	reg v_keyinput_19_v;
	reg v_keyinput_20_v;
	reg v_keyinput_21_v;
	reg v_keyinput_22_v;
	reg v_keyinput_23_v;
	reg v_keyinput_24_v;
	reg v_keyinput_25_v;
	reg v_keyinput_26_v;
	reg v_keyinput_27_v;
	reg v_keyinput_28_v;
	reg v_keyinput_29_v;
	reg v_keyinput_30_v;
	reg v_keyinput_31_v;
	reg v_keyinput_32_v;
	reg v_keyinput_33_v;
	reg v_keyinput_34_v;
	reg v_keyinput_35_v;
	reg v_keyinput_36_v;
	reg v_keyinput_37_v;
	reg v_keyinput_38_v;
	reg v_keyinput_39_v;
	reg v_keyinput_40_v;
	reg v_keyinput_41_v;
	reg v_keyinput_42_v;
	reg v_keyinput_43_v;
	reg v_keyinput_44_v;
	reg v_keyinput_45_v;
	reg v_keyinput_46_v;
	reg v_keyinput_47_v;
	reg v_keyinput_48_v;
	reg v_keyinput_49_v;
	reg v_keyinput_50_v;
	reg v_keyinput_51_v;
	reg v_keyinput_52_v;
	reg v_keyinput_53_v;
	reg v_keyinput_54_v;
	reg v_keyinput_55_v;
	reg v_keyinput_56_v;
	reg v_keyinput_57_v;
	reg v_keyinput_58_v;
	reg v_keyinput_59_v;
	reg v_keyinput_60_v;
	reg v_keyinput_61_v;
	reg v_keyinput_62_v;
	reg v_keyinput_63_v;
	reg v_keyinput_64_v;
	reg v_keyinput_65_v;
	reg v_keyinput_66_v;
	reg v_keyinput_67_v;
	reg v_keyinput_68_v;
	reg v_keyinput_69_v;
	reg v_keyinput_70_v;
	reg v_keyinput_71_v;
	reg v_keyinput_72_v;
	reg v_keyinput_73_v;
	reg v_keyinput_74_v;
	reg v_keyinput_75_v;
	reg v_keyinput_76_v;
	reg v_keyinput_77_v;
	reg v_keyinput_78_v;
	reg v_keyinput_79_v;
	reg v_keyinput_80_v;
	reg v_keyinput_81_v;
	reg v_keyinput_82_v;
	reg v_keyinput_83_v;
	reg v_keyinput_84_v;
	reg v_keyinput_85_v;
	reg v_keyinput_86_v;
	reg v_keyinput_87_v;
	reg v_keyinput_88_v;
	reg v_keyinput_89_v;
	reg v_keyinput_90_v;
	reg v_keyinput_91_v;
	reg v_keyinput_92_v;
	reg v_keyinput_93_v;
	reg v_keyinput_94_v;
	reg v_keyinput_95_v;
	reg v_keyinput_96_v;
	reg v_keyinput_97_v;
	reg v_keyinput_98_v;
	reg v_keyinput_99_v;
	reg v_keyinput_100_v;
	reg v_keyinput_101_v;
	reg v_keyinput_102_v;
	reg v_keyinput_103_v;
	reg v_keyinput_104_v;
	reg v_keyinput_105_v;
	reg v_keyinput_106_v;
	reg v_keyinput_107_v;
	reg v_keyinput_108_v;
	reg v_keyinput_109_v;
	reg v_keyinput_110_v;
	reg v_keyinput_111_v;
	reg v_keyinput_112_v;
	reg v_keyinput_113_v;
	reg v_keyinput_114_v;
	reg v_keyinput_115_v;
	reg v_keyinput_116_v;
	reg v_keyinput_117_v;
	reg v_keyinput_118_v;
	reg v_keyinput_119_v;
	reg v_keyinput_120_v;
	reg v_keyinput_121_v;
	reg v_keyinput_122_v;
	reg v_keyinput_123_v;
	reg v_keyinput_124_v;
	reg v_keyinput_125_v;
	reg v_keyinput_126_v;
	reg v_keyinput_127_v;

  // Outputs
  wire v_o1_v;
	wire v_o2_v;
	wire v_o3_v;
	wire v_o4_v;
	wire v_o5_v;
	wire v_o6_v;
	wire v_o7_v;
	wire v_o8_v;
	wire v_o9_v;
	wire v_o10_v;
	wire v_o11_v;
	wire v_o12_v;
	wire v_o13_v;
	wire v_o14_v;
	wire v_o15_v;
	wire v_o16_v;
	wire v_o17_v;
	wire v_o18_v;
	wire v_o19_v;
	wire v_o20_v;
	wire v_o21_v;
	wire v_o22_v;

  reg [182:0] read_data [0:0];
	integer i;
	integer write_data;

  // Clock and reset signals
  reg v_in1_v;
  reg rst;
  integer file;

  // Instantiate the Design Under Test (DUT)
  circuit_design UUT (
    .reset(rst),
    .v_in1_v(v_in1_v),
    .v_in2_v(v_in2_v), 
    .v_in3_v(v_in3_v), 
    .v_in4_v(v_in4_v), 
    .v_in5_v(v_in5_v), 
    .v_in6_v(v_in6_v), 
    .v_in7_v(v_in7_v), 
    .v_in8_v(v_in8_v), 
    .v_in9_v(v_in9_v), 
    .v_in10_v(v_in10_v), 
    .v_in11_v(v_in11_v), 
    .v_in12_v(v_in12_v), 
    .v_in13_v(v_in13_v), 
    .v_in14_v(v_in14_v), 
    .v_in15_v(v_in15_v), 
    .v_in16_v(v_in16_v), 
    .v_in17_v(v_in17_v), 
    .v_in18_v(v_in18_v), 
    .v_in19_v(v_in19_v), 
    .v_in20_v(v_in20_v), 
    .v_in21_v(v_in21_v), 
    .v_in22_v(v_in22_v), 
    .v_in23_v(v_in23_v), 
    .v_in24_v(v_in24_v), 
    .v_in25_v(v_in25_v), 
    .v_in26_v(v_in26_v), 
    .v_in27_v(v_in27_v), 
    .v_in28_v(v_in28_v), 
    .v_in29_v(v_in29_v), 
    .v_in30_v(v_in30_v), 
    .v_in31_v(v_in31_v), 
    .v_in32_v(v_in32_v), 
    .v_in33_v(v_in33_v), 
    .v_keyinput_0_v(v_keyinput_0_v), 
    .v_keyinput_1_v(v_keyinput_1_v), 
    .v_keyinput_2_v(v_keyinput_2_v), 
    .v_keyinput_3_v(v_keyinput_3_v), 
    .v_keyinput_4_v(v_keyinput_4_v), 
    .v_keyinput_5_v(v_keyinput_5_v), 
    .v_keyinput_6_v(v_keyinput_6_v), 
    .v_keyinput_7_v(v_keyinput_7_v), 
    .v_keyinput_8_v(v_keyinput_8_v), 
    .v_keyinput_9_v(v_keyinput_9_v), 
    .v_keyinput_10_v(v_keyinput_10_v), 
    .v_keyinput_11_v(v_keyinput_11_v), 
    .v_keyinput_12_v(v_keyinput_12_v), 
    .v_keyinput_13_v(v_keyinput_13_v), 
    .v_keyinput_14_v(v_keyinput_14_v), 
    .v_keyinput_15_v(v_keyinput_15_v), 
    .v_keyinput_16_v(v_keyinput_16_v), 
    .v_keyinput_17_v(v_keyinput_17_v), 
    .v_keyinput_18_v(v_keyinput_18_v), 
    .v_keyinput_19_v(v_keyinput_19_v), 
    .v_keyinput_20_v(v_keyinput_20_v), 
    .v_keyinput_21_v(v_keyinput_21_v), 
    .v_keyinput_22_v(v_keyinput_22_v), 
    .v_keyinput_23_v(v_keyinput_23_v), 
    .v_keyinput_24_v(v_keyinput_24_v), 
    .v_keyinput_25_v(v_keyinput_25_v), 
    .v_keyinput_26_v(v_keyinput_26_v), 
    .v_keyinput_27_v(v_keyinput_27_v),
    .v_keyinput_28_v(v_keyinput_28_v),
    .v_keyinput_29_v(v_keyinput_29_v),
    .v_keyinput_30_v(v_keyinput_30_v),
    .v_keyinput_31_v(v_keyinput_31_v),
    .v_keyinput_32_v(v_keyinput_32_v),
    .v_keyinput_33_v(v_keyinput_33_v),
    .v_keyinput_34_v(v_keyinput_34_v),
    .v_keyinput_35_v(v_keyinput_35_v),
    .v_keyinput_36_v(v_keyinput_36_v),
    .v_keyinput_37_v(v_keyinput_37_v),
    .v_keyinput_38_v(v_keyinput_38_v),
    .v_keyinput_39_v(v_keyinput_39_v),
    .v_keyinput_40_v(v_keyinput_40_v),
    .v_keyinput_41_v(v_keyinput_41_v),
    .v_keyinput_42_v(v_keyinput_42_v),
    .v_keyinput_43_v(v_keyinput_43_v),
    .v_keyinput_44_v(v_keyinput_44_v),
    .v_keyinput_45_v(v_keyinput_45_v),
    .v_keyinput_46_v(v_keyinput_46_v),
    .v_keyinput_47_v(v_keyinput_47_v),
    .v_keyinput_48_v(v_keyinput_48_v),
    .v_keyinput_49_v(v_keyinput_49_v),
    .v_keyinput_50_v(v_keyinput_50_v),
    .v_keyinput_51_v(v_keyinput_51_v),
    .v_keyinput_52_v(v_keyinput_52_v),
    .v_keyinput_53_v(v_keyinput_53_v),
    .v_keyinput_54_v(v_keyinput_54_v),
    .v_keyinput_55_v(v_keyinput_55_v),
    .v_keyinput_56_v(v_keyinput_56_v),
    .v_keyinput_57_v(v_keyinput_57_v),
    .v_keyinput_58_v(v_keyinput_58_v),
    .v_keyinput_59_v(v_keyinput_59_v),
    .v_keyinput_60_v(v_keyinput_60_v),
    .v_keyinput_61_v(v_keyinput_61_v),
    .v_keyinput_62_v(v_keyinput_62_v),
    .v_keyinput_63_v(v_keyinput_63_v),
    .v_keyinput_64_v(v_keyinput_64_v),
    .v_keyinput_65_v(v_keyinput_65_v),
    .v_keyinput_66_v(v_keyinput_66_v),
    .v_keyinput_67_v(v_keyinput_67_v),
    .v_keyinput_68_v(v_keyinput_68_v),
    .v_keyinput_69_v(v_keyinput_69_v),
    .v_keyinput_70_v(v_keyinput_70_v),
    .v_keyinput_71_v(v_keyinput_71_v),
    .v_keyinput_72_v(v_keyinput_72_v),
    .v_keyinput_73_v(v_keyinput_73_v),
    .v_keyinput_74_v(v_keyinput_74_v),
    .v_keyinput_75_v(v_keyinput_75_v),
    .v_keyinput_76_v(v_keyinput_76_v),
    .v_keyinput_77_v(v_keyinput_77_v),
    .v_keyinput_78_v(v_keyinput_78_v),
    .v_keyinput_79_v(v_keyinput_79_v),
    .v_keyinput_80_v(v_keyinput_80_v),
    .v_keyinput_81_v(v_keyinput_81_v),
    .v_keyinput_82_v(v_keyinput_82_v),
    .v_keyinput_83_v(v_keyinput_83_v),
    .v_keyinput_84_v(v_keyinput_84_v),
    .v_keyinput_85_v(v_keyinput_85_v),
    .v_keyinput_86_v(v_keyinput_86_v),
    .v_keyinput_87_v(v_keyinput_87_v),
    .v_keyinput_88_v(v_keyinput_88_v),
    .v_keyinput_89_v(v_keyinput_89_v),
    .v_keyinput_90_v(v_keyinput_90_v),
    .v_keyinput_91_v(v_keyinput_91_v),
    .v_keyinput_92_v(v_keyinput_92_v),
    .v_keyinput_93_v(v_keyinput_93_v),
    .v_keyinput_94_v(v_keyinput_94_v),
    .v_keyinput_95_v(v_keyinput_95_v),
    .v_keyinput_96_v(v_keyinput_96_v),
    .v_keyinput_97_v(v_keyinput_97_v),
    .v_keyinput_98_v(v_keyinput_98_v),
    .v_keyinput_99_v(v_keyinput_99_v),
    .v_keyinput_100_v(v_keyinput_100_v),
    .v_keyinput_101_v(v_keyinput_101_v),
    .v_keyinput_102_v(v_keyinput_102_v),
    .v_keyinput_103_v(v_keyinput_103_v),
    .v_keyinput_104_v(v_keyinput_104_v),
    .v_keyinput_105_v(v_keyinput_105_v),
    .v_keyinput_106_v(v_keyinput_106_v),
    .v_keyinput_107_v(v_keyinput_107_v),
    .v_keyinput_108_v(v_keyinput_108_v),
    .v_keyinput_109_v(v_keyinput_109_v),
    .v_keyinput_110_v(v_keyinput_110_v),
    .v_keyinput_111_v(v_keyinput_111_v),
    .v_keyinput_112_v(v_keyinput_112_v),
    .v_keyinput_113_v(v_keyinput_113_v),
    .v_keyinput_114_v(v_keyinput_114_v),
    .v_keyinput_115_v(v_keyinput_115_v),
    .v_keyinput_116_v(v_keyinput_116_v),
    .v_keyinput_117_v(v_keyinput_117_v),
    .v_keyinput_118_v(v_keyinput_118_v),
    .v_keyinput_119_v(v_keyinput_119_v),
    .v_keyinput_120_v(v_keyinput_120_v),
    .v_keyinput_121_v(v_keyinput_121_v),
    .v_keyinput_122_v(v_keyinput_122_v),
    .v_keyinput_123_v(v_keyinput_123_v),
    .v_keyinput_124_v(v_keyinput_124_v),
    .v_keyinput_125_v(v_keyinput_125_v),
    .v_keyinput_126_v(v_keyinput_126_v),
    .v_keyinput_127_v(v_keyinput_127_v),
    .v_o1_v(v_o1_v),
    .v_o2_v(v_o2_v),
    .v_o3_v(v_o3_v),
    .v_o4_v(v_o4_v),
    .v_o5_v(v_o5_v),
    .v_o6_v(v_o6_v),
    .v_o7_v(v_o7_v),
    .v_o8_v(v_o8_v),
    .v_o9_v(v_o9_v),
    .v_o10_v(v_o10_v),
    .v_o11_v(v_o11_v),
    .v_o12_v(v_o12_v),
    .v_o13_v(v_o13_v),
    .v_o14_v(v_o14_v),
    .v_o15_v(v_o15_v),
    .v_o16_v(v_o16_v),
    .v_o17_v(v_o17_v),
    .v_o18_v(v_o18_v),
    .v_o19_v(v_o19_v),
    .v_o20_v(v_o20_v),
    .v_o21_v(v_o21_v),
    .v_o22_v(v_o22_v)
  );

  // Initial values
  initial begin
    $dumpfile("./Execution/large_testBench.vcd");
    $dumpvars(0, testbench);
    file = $fopen("./Execution/large_output.txt", "w");
    v_in1_v = 1;
    $readmemb("./Execution/large_input.txt", read_data);
    { v_in2_v, 
        v_in3_v, 
        v_in4_v, 
        v_in5_v, 
        v_in6_v,
        v_in7_v,
        v_in8_v,
        v_in9_v,
        v_in10_v,
        v_in11_v,
        v_in12_v,
        v_in13_v,
        v_in14_v,
        v_in15_v,
        v_in16_v,
        v_in17_v,
        v_in18_v,
        v_in19_v,
        v_in20_v,
        v_in21_v,
        v_in22_v,
        v_in23_v,
        v_in24_v,
        v_in25_v,
        v_in26_v,
        v_in27_v,
        v_in28_v,
        v_in29_v,
        v_in30_v,
        v_in31_v,
        v_in32_v,
        v_in33_v,
        v_keyinput_0_v,
        v_keyinput_1_v,
        v_keyinput_2_v,
        v_keyinput_3_v,
        v_keyinput_4_v,
        v_keyinput_5_v,
        v_keyinput_6_v,
        v_keyinput_7_v,
        v_keyinput_8_v,
        v_keyinput_9_v,
        v_keyinput_10_v,
        v_keyinput_11_v,
        v_keyinput_12_v,
        v_keyinput_13_v,
        v_keyinput_14_v,
        v_keyinput_15_v,
        v_keyinput_16_v,
        v_keyinput_17_v,
        v_keyinput_18_v,
        v_keyinput_19_v,
        v_keyinput_20_v,
        v_keyinput_21_v,
        v_keyinput_22_v,
        v_keyinput_23_v,
        v_keyinput_24_v,
        v_keyinput_25_v,
        v_keyinput_26_v,
        v_keyinput_27_v,
        v_keyinput_28_v,
        v_keyinput_29_v,
        v_keyinput_30_v,
        v_keyinput_31_v,
        v_keyinput_32_v,
        v_keyinput_33_v,
        v_keyinput_34_v,
        v_keyinput_35_v,
        v_keyinput_36_v,
        v_keyinput_37_v,
        v_keyinput_38_v,
        v_keyinput_39_v,
        v_keyinput_40_v,
        v_keyinput_41_v,
        v_keyinput_42_v,
        v_keyinput_43_v,
        v_keyinput_44_v,
        v_keyinput_45_v,
        v_keyinput_46_v,
        v_keyinput_47_v,
        v_keyinput_48_v,
        v_keyinput_49_v,
        v_keyinput_50_v,
        v_keyinput_51_v,
        v_keyinput_52_v,
        v_keyinput_53_v,
        v_keyinput_54_v,
        v_keyinput_55_v,
        v_keyinput_56_v,
        v_keyinput_57_v,
        v_keyinput_58_v,
        v_keyinput_59_v,
        v_keyinput_60_v,
        v_keyinput_61_v,
        v_keyinput_62_v,
        v_keyinput_63_v,
        v_keyinput_64_v,
        v_keyinput_65_v,
        v_keyinput_66_v,
        v_keyinput_67_v,
        v_keyinput_68_v,
        v_keyinput_69_v,
        v_keyinput_70_v,
        v_keyinput_71_v,
        v_keyinput_72_v,
        v_keyinput_73_v,
        v_keyinput_74_v,
        v_keyinput_75_v,
        v_keyinput_76_v,
        v_keyinput_77_v,
        v_keyinput_78_v,
        v_keyinput_79_v,
        v_keyinput_80_v,
        v_keyinput_81_v,
        v_keyinput_82_v,
        v_keyinput_83_v,
        v_keyinput_84_v,
        v_keyinput_85_v,
        v_keyinput_86_v,
        v_keyinput_87_v,
        v_keyinput_88_v,
        v_keyinput_89_v,
        v_keyinput_90_v,
        v_keyinput_91_v,
        v_keyinput_92_v,
        v_keyinput_93_v,
        v_keyinput_94_v,
        v_keyinput_95_v,
        v_keyinput_96_v,
        v_keyinput_97_v,
        v_keyinput_98_v,
        v_keyinput_99_v,
        v_keyinput_100_v,
        v_keyinput_101_v,
        v_keyinput_102_v,
        v_keyinput_103_v,
        v_keyinput_104_v,
        v_keyinput_105_v,
        v_keyinput_106_v,
        v_keyinput_107_v,
        v_keyinput_108_v,
        v_keyinput_109_v,
        v_keyinput_110_v,
        v_keyinput_111_v,
        v_keyinput_112_v,
        v_keyinput_113_v,
        v_keyinput_114_v,
        v_keyinput_115_v,
        v_keyinput_116_v,
        v_keyinput_117_v,
        v_keyinput_118_v,
        v_keyinput_119_v,
        v_keyinput_120_v,
        v_keyinput_121_v,
        v_keyinput_122_v,
        v_keyinput_123_v,
        v_keyinput_124_v,
        v_keyinput_125_v,
        v_keyinput_126_v,
        v_keyinput_127_v
      } = read_data[0];
    rst = 1;
    #20;
    rst = 0;
  end

  // Clock generator
  always #10 v_in1_v = ~v_in1_v;

  // Test sequence
  always @(posedge v_in1_v) begin
      $fwrite(file, "%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b\n", v_o1_v, v_o2_v, v_o3_v, v_o4_v, v_o5_v, v_o6_v, v_o7_v, v_o8_v, v_o9_v, v_o10_v, v_o11_v, v_o12_v, v_o13_v, v_o14_v, v_o15_v, v_o16_v, v_o17_v, v_o18_v, v_o19_v, v_o20_v, v_o21_v, v_o22_v);
  end 

  initial begin
     #100 
     $fwrite(file, "%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b%b\n", v_o1_v, v_o2_v, v_o3_v, v_o4_v, v_o5_v, v_o6_v, v_o7_v, v_o8_v, v_o9_v, v_o10_v, v_o11_v, v_o12_v, v_o13_v, v_o14_v, v_o15_v, v_o16_v, v_o17_v, v_o18_v, v_o19_v, v_o20_v, v_o21_v, v_o22_v);
     $fclose(file);
     $finish;
  end
endmodule
