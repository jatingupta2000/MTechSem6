`timescale 1ns/10ps//time-unit = 1 ns and precision = 10 ps

module circuit_design(reset, v_in1_v, v_in2_v, v_in3_v, v_in4_v, v_in5_v, v_in6_v, v_in7_v, v_in8_v, v_in9_v, v_in10_v, v_in11_v, v_in12_v, v_in13_v, v_in14_v, v_in15_v, v_in16_v, v_in17_v, v_in18_v, v_in19_v, v_in20_v, v_in21_v, v_in22_v, v_in23_v, v_in24_v, v_in25_v, v_in26_v, v_in27_v, v_in28_v, v_in29_v, v_in30_v, v_in31_v, v_in32_v, v_in33_v, v_keyinput_0_v, v_keyinput_1_v, v_keyinput_2_v, v_keyinput_3_v, v_keyinput_4_v, v_keyinput_5_v, v_keyinput_6_v, v_keyinput_7_v, v_keyinput_8_v, v_keyinput_9_v, v_keyinput_10_v, v_keyinput_11_v, v_keyinput_12_v, v_keyinput_13_v, v_keyinput_14_v, v_keyinput_15_v, v_keyinput_16_v, v_keyinput_17_v, v_keyinput_18_v, v_keyinput_19_v, v_keyinput_20_v, v_keyinput_21_v, v_keyinput_22_v, v_keyinput_23_v, v_keyinput_24_v, v_keyinput_25_v, v_keyinput_26_v, v_keyinput_27_v, v_keyinput_28_v, v_keyinput_29_v, v_keyinput_30_v, v_keyinput_31_v, v_keyinput_32_v, v_keyinput_33_v, v_keyinput_34_v, v_keyinput_35_v, v_keyinput_36_v, v_keyinput_37_v, v_keyinput_38_v, v_keyinput_39_v, v_keyinput_40_v, v_keyinput_41_v, v_keyinput_42_v, v_keyinput_43_v, v_keyinput_44_v, v_keyinput_45_v, v_keyinput_46_v, v_keyinput_47_v, v_keyinput_48_v, v_keyinput_49_v, v_keyinput_50_v, v_keyinput_51_v, v_keyinput_52_v, v_keyinput_53_v, v_keyinput_54_v, v_keyinput_55_v, v_keyinput_56_v, v_keyinput_57_v, v_keyinput_58_v, v_keyinput_59_v, v_keyinput_60_v, v_keyinput_61_v, v_keyinput_62_v, v_keyinput_63_v, v_keyinput_64_v, v_keyinput_65_v, v_keyinput_66_v, v_keyinput_67_v, v_keyinput_68_v, v_keyinput_69_v, v_keyinput_70_v, v_keyinput_71_v, v_keyinput_72_v, v_keyinput_73_v, v_keyinput_74_v, v_keyinput_75_v, v_keyinput_76_v, v_keyinput_77_v, v_keyinput_78_v, v_keyinput_79_v, v_keyinput_80_v, v_keyinput_81_v, v_keyinput_82_v, v_keyinput_83_v, v_keyinput_84_v, v_keyinput_85_v, v_keyinput_86_v, v_keyinput_87_v, v_keyinput_88_v, v_keyinput_89_v, v_keyinput_90_v, v_keyinput_91_v, v_keyinput_92_v, v_keyinput_93_v, v_keyinput_94_v, v_keyinput_95_v, v_keyinput_96_v, v_keyinput_97_v, v_keyinput_98_v, v_keyinput_99_v, v_keyinput_100_v, v_keyinput_101_v, v_keyinput_102_v, v_keyinput_103_v, v_keyinput_104_v, v_keyinput_105_v, v_keyinput_106_v, v_keyinput_107_v, v_keyinput_108_v, v_keyinput_109_v, v_keyinput_110_v, v_keyinput_111_v, v_keyinput_112_v, v_keyinput_113_v, v_keyinput_114_v, v_keyinput_115_v, v_keyinput_116_v, v_keyinput_117_v, v_keyinput_118_v, v_keyinput_119_v, v_keyinput_120_v, v_keyinput_121_v, v_keyinput_122_v, v_keyinput_123_v, v_keyinput_124_v, v_keyinput_125_v, v_keyinput_126_v, v_keyinput_127_v, v_o1_v, v_o2_v, v_o3_v, v_o4_v, v_o5_v, v_o6_v, v_o7_v, v_o8_v, v_o9_v, v_o10_v, v_o11_v, v_o12_v, v_o13_v, v_o14_v, v_o15_v, v_o16_v, v_o17_v, v_o18_v, v_o19_v, v_o20_v, v_o21_v, v_o22_v);
	input reset;
	input v_in1_v;
	input v_in2_v;
	input v_in3_v;
	input v_in4_v;
	input v_in5_v;
	input v_in6_v;
	input v_in7_v;
	input v_in8_v;
	input v_in9_v;
	input v_in10_v;
	input v_in11_v;
	input v_in12_v;
	input v_in13_v;
	input v_in14_v;
	input v_in15_v;
	input v_in16_v;
	input v_in17_v;
	input v_in18_v;
	input v_in19_v;
	input v_in20_v;
	input v_in21_v;
	input v_in22_v;
	input v_in23_v;
	input v_in24_v;
	input v_in25_v;
	input v_in26_v;
	input v_in27_v;
	input v_in28_v;
	input v_in29_v;
	input v_in30_v;
	input v_in31_v;
	input v_in32_v;
	input v_in33_v;
	input v_keyinput_0_v;
	input v_keyinput_1_v;
	input v_keyinput_2_v;
	input v_keyinput_3_v;
	input v_keyinput_4_v;
	input v_keyinput_5_v;
	input v_keyinput_6_v;
	input v_keyinput_7_v;
	input v_keyinput_8_v;
	input v_keyinput_9_v;
	input v_keyinput_10_v;
	input v_keyinput_11_v;
	input v_keyinput_12_v;
	input v_keyinput_13_v;
	input v_keyinput_14_v;
	input v_keyinput_15_v;
	input v_keyinput_16_v;
	input v_keyinput_17_v;
	input v_keyinput_18_v;
	input v_keyinput_19_v;
	input v_keyinput_20_v;
	input v_keyinput_21_v;
	input v_keyinput_22_v;
	input v_keyinput_23_v;
	input v_keyinput_24_v;
	input v_keyinput_25_v;
	input v_keyinput_26_v;
	input v_keyinput_27_v;
	input v_keyinput_28_v;
	input v_keyinput_29_v;
	input v_keyinput_30_v;
	input v_keyinput_31_v;
	input v_keyinput_32_v;
	input v_keyinput_33_v;
	input v_keyinput_34_v;
	input v_keyinput_35_v;
	input v_keyinput_36_v;
	input v_keyinput_37_v;
	input v_keyinput_38_v;
	input v_keyinput_39_v;
	input v_keyinput_40_v;
	input v_keyinput_41_v;
	input v_keyinput_42_v;
	input v_keyinput_43_v;
	input v_keyinput_44_v;
	input v_keyinput_45_v;
	input v_keyinput_46_v;
	input v_keyinput_47_v;
	input v_keyinput_48_v;
	input v_keyinput_49_v;
	input v_keyinput_50_v;
	input v_keyinput_51_v;
	input v_keyinput_52_v;
	input v_keyinput_53_v;
	input v_keyinput_54_v;
	input v_keyinput_55_v;
	input v_keyinput_56_v;
	input v_keyinput_57_v;
	input v_keyinput_58_v;
	input v_keyinput_59_v;
	input v_keyinput_60_v;
	input v_keyinput_61_v;
	input v_keyinput_62_v;
	input v_keyinput_63_v;
	input v_keyinput_64_v;
	input v_keyinput_65_v;
	input v_keyinput_66_v;
	input v_keyinput_67_v;
	input v_keyinput_68_v;
	input v_keyinput_69_v;
	input v_keyinput_70_v;
	input v_keyinput_71_v;
	input v_keyinput_72_v;
	input v_keyinput_73_v;
	input v_keyinput_74_v;
	input v_keyinput_75_v;
	input v_keyinput_76_v;
	input v_keyinput_77_v;
	input v_keyinput_78_v;
	input v_keyinput_79_v;
	input v_keyinput_80_v;
	input v_keyinput_81_v;
	input v_keyinput_82_v;
	input v_keyinput_83_v;
	input v_keyinput_84_v;
	input v_keyinput_85_v;
	input v_keyinput_86_v;
	input v_keyinput_87_v;
	input v_keyinput_88_v;
	input v_keyinput_89_v;
	input v_keyinput_90_v;
	input v_keyinput_91_v;
	input v_keyinput_92_v;
	input v_keyinput_93_v;
	input v_keyinput_94_v;
	input v_keyinput_95_v;
	input v_keyinput_96_v;
	input v_keyinput_97_v;
	input v_keyinput_98_v;
	input v_keyinput_99_v;
	input v_keyinput_100_v;
	input v_keyinput_101_v;
	input v_keyinput_102_v;
	input v_keyinput_103_v;
	input v_keyinput_104_v;
	input v_keyinput_105_v;
	input v_keyinput_106_v;
	input v_keyinput_107_v;
	input v_keyinput_108_v;
	input v_keyinput_109_v;
	input v_keyinput_110_v;
	input v_keyinput_111_v;
	input v_keyinput_112_v;
	input v_keyinput_113_v;
	input v_keyinput_114_v;
	input v_keyinput_115_v;
	input v_keyinput_116_v;
	input v_keyinput_117_v;
	input v_keyinput_118_v;
	input v_keyinput_119_v;
	input v_keyinput_120_v;
	input v_keyinput_121_v;
	input v_keyinput_122_v;
	input v_keyinput_123_v;
	input v_keyinput_124_v;
	input v_keyinput_125_v;
	input v_keyinput_126_v;
	input v_keyinput_127_v;
	output v_o1_v;
	output v_o2_v;
	output v_o3_v;
	output v_o4_v;
	output v_o5_v;
	output v_o6_v;
	output v_o7_v;
	output v_o8_v;
	output v_o9_v;
	output v_o10_v;
	output v_o11_v;
	output v_o12_v;
	output v_o13_v;
	output v_o14_v;
	output v_o15_v;
	output v_o16_v;
	output v_o17_v;
	output v_o18_v;
	output v_o19_v;
	output v_o20_v;
	output v_o21_v;
	output v_o22_v;
	wire v_w6528_v;
	wire v_w5688_v;
	wire v_w1019_v;
	wire v_w4890_v;
	wire v_w3972_v;
	wire v_w7621_v;
	wire v_w7678_v;
	wire v_w6429_v;
	wire v_w814_v;
	wire v_w6766_v;
	wire v_w7341_v;
	wire v_w5016_v;
	wire v_w3944_v;
	wire v_w4594_v;
	wire v_w5353_v;
	wire v_w1417_v;
	wire v_w2068_v;
	wire v_w7007_v;
	wire v_w4360_v;
	wire v_w1888_v;
	reg v_s263_v;
	wire v_w3434_v;
	wire v_w1243_v;
	wire v_w1519_v;
	wire v_w6954_v;
	wire v_w6248_v;
	wire v_w8086_v;
	wire v_w1296_v;
	wire v_w4224_v;
	wire v_w7289_v;
	wire v_w6507_v;
	wire v_w314_v;
	wire v_w4236_v;
	wire v_w7834_v;
	wire v_w6135_v;
	wire v_w6143_v;
	wire v_w5844_v;
	wire v_w2771_v;
	wire v_w3120_v;
	wire v_w5487_v;
	wire v_w5965_v;
	wire v_w445_v;
	wire v_w7554_v;
	wire v_w1688_v;
	wire v_w3768_v;
	wire v_w8160_v;
	wire v_w8229_v;
	wire v_w4354_v;
	wire v_w2930_v;
	wire v_w5471_v;
	wire v_w2154_v;
	wire v_w121_v;
	wire v_w3505_v;
	wire v_w5873_v;
	wire v_w7027_v;
	wire v_w7211_v;
	wire v_w2600_v;
	wire v_w6819_v;
	wire v_w6346_v;
	wire v_w1290_v;
	wire v_w3979_v;
	wire v_w2244_v;
	wire v_w7366_v;
	wire v_w5477_v;
	wire v_w6103_v;
	reg v_s19_v;
	reg v_s39_v;
	wire v_w4834_v;
	wire v_w3523_v;
	wire v_w7525_v;
	wire v_w708_v;
	wire v_w5945_v;
	wire v_w442_v;
	reg v_s455_v;
	wire v_w5609_v;
	wire v_w4734_v;
	wire v_w7244_v;
	wire v_w1740_v;
	wire v_w794_v;
	wire v_w7374_v;
	wire v_w6797_v;
	wire v_w643_v;
	wire v_w7229_v;
	wire v_w5578_v;
	wire v_w2127_v;
	wire v_w2296_v;
	wire v_w4635_v;
	wire v_w1733_v;
	wire v_w3456_v;
	wire v_w1552_v;
	wire v_w7474_v;
	wire v_w5762_v;
	wire v_w1883_v;
	wire v_w4446_v;
	wire v_w2471_v;
	wire v_w450_v;
	wire v_w6544_v;
	wire v_w2176_v;
	wire v_w6105_v;
	wire v_w6756_v;
	wire v_w612_v;
	wire v_w4157_v;
	wire v_w429_v;
	wire v_w3415_v;
	wire v_w1122_v;
	wire v_w5283_v;
	wire v_w2926_v;
	wire v_w1823_v;
	wire v_w551_v;
	reg v_s488_v;
	wire v_w3073_v;
	wire v_w8222_v;
	wire v_w3152_v;
	wire v_w308_v;
	wire v_w4670_v;
	wire v_w5865_v;
	wire v_w5784_v;
	wire v_w7556_v;
	wire v_w2378_v;
	wire v_w7097_v;
	reg v_s456_v;
	wire v_w3180_v;
	wire v_w3620_v;
	wire v_w7240_v;
	wire v_w2259_v;
	wire v_w5582_v;
	wire v_w5871_v;
	wire v_w6695_v;
	wire v_w628_v;
	wire v_w4772_v;
	wire v_w7989_v;
	wire v_w8178_v;
	wire v_w8159_v;
	wire v_w1371_v;
	wire v_w2763_v;
	wire v_w6527_v;
	wire v_w947_v;
	wire v_w5932_v;
	wire v_w5731_v;
	wire v_w6674_v;
	wire v_w3286_v;
	wire v_w224_v;
	wire v_w3255_v;
	wire v_w7472_v;
	wire v_w5170_v;
	wire v_w4709_v;
	wire v_w4866_v;
	wire v_w6564_v;
	wire v_w6316_v;
	wire v_w2518_v;
	wire v_w3722_v;
	wire v_w1884_v;
	wire v_w6147_v;
	wire v_w1024_v;
	wire v_w6524_v;
	wire v_w2352_v;
	wire v_w1175_v;
	wire v_w7662_v;
	wire v_w3994_v;
	wire v_w8028_v;
	wire v_w681_v;
	wire v_w1030_v;
	wire v_w1693_v;
	wire v_w3197_v;
	wire v_w1113_v;
	wire v_w5661_v;
	wire v_w7266_v;
	wire v_w3269_v;
	wire v_w4180_v;
	wire v_w6946_v;
	wire v_w7043_v;
	wire v_w3715_v;
	wire v_w4388_v;
	wire v_w3587_v;
	wire v_w463_v;
	wire v_w4712_v;
	wire v_w3922_v;
	wire v_w5842_v;
	wire v_w2356_v;
	wire v_w1634_v;
	wire v_w607_v;
	wire v_w7731_v;
	wire v_w425_v;
	wire v_w7416_v;
	wire v_w6120_v;
	wire v_w3013_v;
	wire v_w2325_v;
	wire v_w2819_v;
	wire v_w5937_v;
	wire v_w1559_v;
	wire v_w1315_v;
	wire v_w5763_v;
	wire v_w3877_v;
	wire v_w35_v;
	wire v_w3309_v;
	wire v_w2770_v;
	wire v_w1053_v;
	wire v_w6436_v;
	wire v_w3435_v;
	wire v_w6432_v;
	wire v_w3099_v;
	wire v_w5713_v;
	wire v_w5252_v;
	wire v_w3955_v;
	reg v_s45_v;
	reg v_s8_v;
	wire v_w2245_v;
	wire v_w648_v;
	wire v_w4165_v;
	wire v_w1202_v;
	wire v_w1485_v;
	wire v_w6475_v;
	wire v_w1587_v;
	wire v_w4675_v;
	wire v_w5654_v;
	wire v_w7938_v;
	wire v_w3335_v;
	wire v_w1165_v;
	wire v_w6042_v;
	wire v_w705_v;
	wire v_w3832_v;
	wire v_w4320_v;
	wire v_w3028_v;
	wire v_w6688_v;
	wire v_w2338_v;
	wire v_w6447_v;
	wire v_w7033_v;
	wire v_w5900_v;
	wire v_w6362_v;
	reg v_s512_v;
	wire v_w2517_v;
	wire v_w3017_v;
	wire v_w2659_v;
	wire v_w3607_v;
	wire v_w3990_v;
	wire v_w7055_v;
	wire v_w4074_v;
	wire v_w1919_v;
	wire v_w6405_v;
	wire v_w227_v;
	wire v_w2519_v;
	wire v_w2668_v;
	wire v_w1725_v;
	reg v_s273_v;
	wire v_w6372_v;
	wire v_w4751_v;
	wire v_w6560_v;
	wire v_w1676_v;
	wire v_w2617_v;
	wire v_w2532_v;
	wire v_w3401_v;
	wire v_w3347_v;
	wire v_w4099_v;
	wire v_w4854_v;
	wire v_w5437_v;
	reg v_s124_v;
	wire v_w5410_v;
	wire v_w2308_v;
	wire v_w3399_v;
	wire v_w5878_v;
	wire v_w1082_v;
	wire v_w2415_v;
	wire v_w6577_v;
	wire v_w1263_v;
	wire v_w5478_v;
	wire v_w6400_v;
	wire v_w2753_v;
	wire v_w2558_v;
	wire v_w4049_v;
	wire v_w7287_v;
	reg v_s449_v;
	wire v_w2345_v;
	wire v_w5129_v;
	wire v_w5012_v;
	reg v_s94_v;
	wire v_w1821_v;
	wire v_w454_v;
	wire v_w4747_v;
	wire v_w7003_v;
	reg v_s374_v;
	wire v_w6461_v;
	wire v_w3561_v;
	wire v_w2290_v;
	wire v_w6733_v;
	wire v_w8087_v;
	wire v_w4065_v;
	wire v_w4192_v;
	wire v_w5628_v;
	wire v_w7483_v;
	wire v_w7471_v;
	wire v_w1624_v;
	wire v_w3361_v;
	wire v_w3353_v;
	wire v_w2094_v;
	wire v_w2703_v;
	wire v_w4036_v;
	wire v_w5860_v;
	wire v_w3894_v;
	wire v_w1851_v;
	wire v_w4400_v;
	wire v_w4061_v;
	wire v_w1869_v;
	wire v_w3215_v;
	reg v_s511_v;
	wire v_w7870_v;
	wire v_w4417_v;
	wire v_w2886_v;
	wire v_w5841_v;
	wire v_w241_v;
	wire v_w2293_v;
	wire v_w2485_v;
	wire v_w6171_v;
	wire v_w3754_v;
	wire v_w6011_v;
	wire v_w8174_v;
	wire v_w5585_v;
	wire v_w7915_v;
	wire v_w8079_v;
	wire v_w48_v;
	wire v_w5852_v;
	wire v_w2097_v;
	wire v_w3619_v;
	wire v_w2339_v;
	wire v_w4889_v;
	wire v_w8197_v;
	reg v_s65_v;
	wire v_w4468_v;
	wire v_w1592_v;
	wire v_w6419_v;
	wire v_w4525_v;
	wire v_w769_v;
	wire v_w1595_v;
	wire v_w8151_v;
	wire v_w5599_v;
	wire v_w4155_v;
	wire v_w600_v;
	wire v_w6045_v;
	wire v_w7458_v;
	wire v_w3723_v;
	reg v_s43_v;
	wire v_w5926_v;
	wire v_w6251_v;
	wire v_w1757_v;
	wire v_w2088_v;
	wire v_w6304_v;
	wire v_w5118_v;
	wire v_w1801_v;
	wire v_w3189_v;
	wire v_w322_v;
	wire v_w1984_v;
	wire v_w7926_v;
	wire v_w7701_v;
	wire v_w2228_v;
	wire v_w2714_v;
	wire v_w3991_v;
	reg v_s35_v;
	wire v_w3314_v;
	wire v_w397_v;
	wire v_w7037_v;
	wire v_w6683_v;
	wire v_w7503_v;
	wire v_w5491_v;
	wire v_w5619_v;
	wire v_w7986_v;
	reg v_s229_v;
	wire v_w4754_v;
	wire v_w2041_v;
	wire v_w4330_v;
	wire v_w7572_v;
	wire v_w6569_v;
	wire v_w878_v;
	wire v_w882_v;
	wire v_w391_v;
	wire v_w4685_v;
	wire v_w5825_v;
	wire v_w3018_v;
	wire v_w2089_v;
	wire v_w4644_v;
	wire v_w3733_v;
	wire v_w496_v;
	wire v_w6791_v;
	reg v_s238_v;
	wire v_w3240_v;
	wire v_w4498_v;
	wire v_w6210_v;
	wire v_w2144_v;
	wire v_w4613_v;
	wire v_w2492_v;
	wire v_w7052_v;
	wire v_w5698_v;
	wire v_w3397_v;
	wire v_w2759_v;
	wire v_w3293_v;
	wire v_w3104_v;
	reg v_s402_v;
	wire v_w4237_v;
	wire v_w7590_v;
	wire v_w4208_v;
	wire v_w3662_v;
	wire v_w2723_v;
	wire v_w6130_v;
	wire v_w6058_v;
	wire v_w4177_v;
	wire v_w3468_v;
	wire v_w5242_v;
	wire v_w928_v;
	reg v_s308_v;
	wire v_w8071_v;
	wire v_w3525_v;
	wire v_w7610_v;
	wire v_w4748_v;
	reg v_s29_v;
	wire v_w216_v;
	wire v_w618_v;
	wire v_w5635_v;
	wire v_w1542_v;
	wire v_w2929_v;
	wire v_w4797_v;
	wire v_w6862_v;
	wire v_w332_v;
	wire v_w6299_v;
	wire v_w1640_v;
	reg v_s160_v;
	reg v_s78_v;
	wire v_w3362_v;
	wire v_w2712_v;
	wire v_w7467_v;
	wire v_w961_v;
	reg v_s48_v;
	wire v_w3040_v;
	wire v_w6639_v;
	wire v_w7798_v;
	wire v_w4173_v;
	wire v_w6074_v;
	wire v_w6197_v;
	wire v_w5553_v;
	wire v_w5150_v;
	reg v_s165_v;
	wire v_w344_v;
	wire v_w5790_v;
	wire v_w6580_v;
	wire v_w1357_v;
	wire v_w1925_v;
	wire v_w630_v;
	wire v_w3650_v;
	wire v_w240_v;
	wire v_w2900_v;
	wire v_w7772_v;
	wire v_w1711_v;
	wire v_w8111_v;
	wire v_w8194_v;
	wire v_w7505_v;
	wire v_w3524_v;
	wire v_w2936_v;
	wire v_w3985_v;
	wire v_w7825_v;
	wire v_w6458_v;
	wire v_w1306_v;
	wire v_w4136_v;
	wire v_w6153_v;
	wire v_w2794_v;
	wire v_w428_v;
	wire v_w6076_v;
	wire v_w5779_v;
	wire v_w1989_v;
	wire v_w3109_v;
	wire v_w5758_v;
	wire v_w1950_v;
	wire v_w7905_v;
	wire v_w5320_v;
	wire v_w8014_v;
	wire v_w5803_v;
	wire v_w1755_v;
	wire v_w5969_v;
	wire v_w7405_v;
	wire v_w3491_v;
	wire v_w8055_v;
	reg v_s445_v;
	wire v_w5962_v;
	wire v_w4930_v;
	wire v_w4682_v;
	reg v_s409_v;
	wire v_w3012_v;
	wire v_w6525_v;
	wire v_w3960_v;
	wire v_w3190_v;
	wire v_w4238_v;
	reg v_s231_v;
	wire v_w1739_v;
	reg v_s144_v;
	wire v_w7614_v;
	wire v_w8210_v;
	wire v_w4634_v;
	wire v_w7671_v;
	wire v_w4698_v;
	wire v_w672_v;
	wire v_w6053_v;
	wire v_w2316_v;
	wire v_w5017_v;
	wire v_w1828_v;
	wire v_w7491_v;
	wire v_w840_v;
	wire v_w3829_v;
	wire v_w2957_v;
	wire v_w7673_v;
	wire v_w3171_v;
	wire v_w7428_v;
	wire v_w5830_v;
	wire v_w6082_v;
	wire v_w6691_v;
	wire v_w30_v;
	wire v_w5375_v;
	wire v_w2962_v;
	wire v_w1073_v;
	wire v_w4046_v;
	reg v_s351_v;
	wire v_w103_v;
	wire v_w441_v;
	wire v_w3093_v;
	wire v_w7169_v;
	wire v_w5704_v;
	wire v_w7132_v;
	wire v_w6063_v;
	wire v_w2526_v;
	reg v_s138_v;
	wire v_w587_v;
	wire v_w1460_v;
	wire v_w8204_v;
	reg v_s339_v;
	wire v_w1562_v;
	wire v_w1710_v;
	wire v_w3676_v;
	wire v_w5259_v;
	wire v_w2482_v;
	wire v_w1896_v;
	wire v_w1853_v;
	wire v_w1043_v;
	wire v_w3264_v;
	wire v_w3043_v;
	wire v_w1379_v;
	wire v_w8039_v;
	reg v_s122_v;
	wire v_w3632_v;
	wire v_w4019_v;
	wire v_w8135_v;
	wire v_w5389_v;
	wire v_w1117_v;
	wire v_w4279_v;
	wire v_w4804_v;
	wire v_w2387_v;
	wire v_w305_v;
	wire v_w7304_v;
	wire v_w5106_v;
	wire v_w265_v;
	wire v_w1759_v;
	wire v_w1897_v;
	wire v_w6264_v;
	reg v_s434_v;
	wire v_w5961_v;
	reg v_s83_v;
	wire v_w2541_v;
	reg v_s267_v;
	wire v_w8184_v;
	wire v_w4084_v;
	reg v_s173_v;
	wire v_w6654_v;
	wire v_w2530_v;
	wire v_w3720_v;
	wire v_w1861_v;
	wire v_w7773_v;
	wire v_w7080_v;
	wire v_w5429_v;
	wire v_w507_v;
	wire v_w7606_v;
	wire v_w5870_v;
	wire v_w6136_v;
	wire v_w1966_v;
	wire v_w1333_v;
	wire v_w5450_v;
	wire v_w175_v;
	wire v_w1129_v;
	wire v_w6094_v;
	wire v_w60_v;
	wire v_w3901_v;
	wire v_w7456_v;
	wire v_w903_v;
	wire v_w3233_v;
	wire v_w6485_v;
	wire v_w475_v;
	wire v_w4287_v;
	wire v_w7839_v;
	wire v_w4458_v;
	wire v_w5356_v;
	wire v_w874_v;
	wire v_w4473_v;
	wire v_w3648_v;
	wire v_w3500_v;
	wire v_w4620_v;
	wire v_w3970_v;
	wire v_w6649_v;
	wire v_w7794_v;
	wire v_w6018_v;
	reg v_s219_v;
	wire v_w1131_v;
	wire v_w7306_v;
	wire v_w5203_v;
	wire v_w2878_v;
	wire v_w1097_v;
	wire v_w7913_v;
	wire v_w6520_v;
	wire v_w7410_v;
	wire v_w62_v;
	reg v_s400_v;
	wire v_w1526_v;
	wire v_w3695_v;
	wire v_w8069_v;
	wire v_w5883_v;
	wire v_w4048_v;
	wire v_w5594_v;
	wire v_w8148_v;
	wire v_w761_v;
	wire v_w8219_v;
	wire v_w4971_v;
	wire v_w3466_v;
	wire v_w2187_v;
	wire v_w6543_v;
	wire v_w2038_v;
	wire v_w3089_v;
	wire v_w2112_v;
	wire v_w5004_v;
	wire v_w7162_v;
	wire v_w2263_v;
	wire v_w6774_v;
	wire v_w3625_v;
	wire v_w7264_v;
	wire v_w788_v;
	wire v_w983_v;
	wire v_w7478_v;
	wire v_w2233_v;
	wire v_w4875_v;
	wire v_w4103_v;
	wire v_w3129_v;
	wire v_w1191_v;
	wire v_w3674_v;
	wire v_w323_v;
	wire v_w7143_v;
	wire v_w2285_v;
	wire v_w6771_v;
	wire v_w6588_v;
	wire v_w512_v;
	wire v_w3003_v;
	wire v_w2594_v;
	wire v_w5197_v;
	wire v_w5226_v;
	wire v_w189_v;
	wire v_w8120_v;
	wire v_w1160_v;
	wire v_w1997_v;
	wire v_w5580_v;
	wire v_w5430_v;
	wire v_w4247_v;
	wire v_w2484_v;
	wire v_w1647_v;
	wire v_w5753_v;
	wire v_w7804_v;
	wire v_w1092_v;
	wire v_w1572_v;
	wire v_w4835_v;
	wire v_w8179_v;
	wire v_w3462_v;
	wire v_w5575_v;
	wire v_w3363_v;
	wire v_w4781_v;
	wire v_w2809_v;
	reg v_s426_v;
	wire v_w2490_v;
	wire v_w3409_v;
	wire v_w2267_v;
	wire v_w5318_v;
	wire v_w1837_v;
	wire v_w4555_v;
	wire v_w6979_v;
	wire v_w2209_v;
	wire v_w5563_v;
	wire v_w201_v;
	wire v_w7021_v;
	wire v_w7544_v;
	wire v_w7685_v;
	wire v_w7068_v;
	wire v_w7784_v;
	wire v_w1013_v;
	wire v_w2065_v;
	wire v_w2194_v;
	wire v_w653_v;
	reg v_s296_v;
	wire v_w6832_v;
	wire v_w6282_v;
	wire v_w285_v;
	wire v_w2095_v;
	wire v_w1909_v;
	wire v_w1496_v;
	wire v_w6384_v;
	wire v_w1674_v;
	wire v_w5548_v;
	wire v_w5497_v;
	wire v_w4430_v;
	wire v_w2707_v;
	wire v_w4575_v;
	wire v_w7220_v;
	wire v_w4438_v;
	wire v_w5928_v;
	wire v_w1846_v;
	wire v_w6966_v;
	wire v_w6775_v;
	wire v_w2320_v;
	reg v_s217_v;
	wire v_w3567_v;
	wire v_w6027_v;
	wire v_w4809_v;
	wire v_w6534_v;
	wire v_w7812_v;
	wire v_w4970_v;
	wire v_w4367_v;
	wire v_w1528_v;
	wire v_w4396_v;
	wire v_w4393_v;
	wire v_w166_v;
	wire v_w6487_v;
	wire v_w1232_v;
	wire v_w1023_v;
	wire v_w7050_v;
	wire v_w2953_v;
	wire v_w4130_v;
	wire v_w2303_v;
	wire v_w1800_v;
	wire v_w3298_v;
	wire v_w273_v;
	wire v_w3137_v;
	wire v_w5273_v;
	wire v_w1108_v;
	wire v_w6486_v;
	wire v_w4187_v;
	wire v_w1394_v;
	wire v_w7020_v;
	wire v_w6730_v;
	wire v_w5571_v;
	wire v_w7342_v;
	wire v_w7029_v;
	reg v_s429_v;
	wire v_w3176_v;
	reg v_s59_v;
	wire v_w5394_v;
	wire v_w7517_v;
	wire v_w2963_v;
	wire v_w730_v;
	wire v_w3791_v;
	wire v_w5804_v;
	wire v_w5902_v;
	wire v_w7843_v;
	wire v_w4045_v;
	wire v_w7243_v;
	wire v_w4795_v;
	wire v_w583_v;
	wire v_w3404_v;
	wire v_w1398_v;
	wire v_w1432_v;
	wire v_w1464_v;
	wire v_w7072_v;
	reg v_s320_v;
	wire v_w6000_v;
	wire v_w7088_v;
	wire v_w5298_v;
	wire v_w6653_v;
	wire v_w1436_v;
	wire v_w2092_v;
	wire v_w7751_v;
	wire v_w857_v;
	wire v_w2029_v;
	wire v_w3250_v;
	wire v_w2146_v;
	wire v_w7446_v;
	wire v_w6944_v;
	wire v_w7880_v;
	wire v_w3421_v;
	wire v_w2162_v;
	wire v_w6650_v;
	wire v_w3705_v;
	wire v_w6266_v;
	wire v_w4090_v;
	wire v_w145_v;
	wire v_w2108_v;
	wire v_w2499_v;
	wire v_w654_v;
	wire v_w6915_v;
	wire v_w6682_v;
	wire v_w3273_v;
	wire v_w6491_v;
	wire v_w6921_v;
	wire v_w8091_v;
	wire v_w5238_v;
	wire v_w7395_v;
	wire v_w8164_v;
	wire v_w2645_v;
	wire v_w2789_v;
	wire v_w110_v;
	wire v_w7699_v;
	wire v_w3126_v;
	wire v_w2540_v;
	wire v_w1876_v;
	wire v_w5561_v;
	wire v_w6790_v;
	wire v_w251_v;
	wire v_w4691_v;
	wire v_w3666_v;
	wire v_w5985_v;
	wire v_w5365_v;
	wire v_w6012_v;
	wire v_w3967_v;
	wire v_w4792_v;
	wire v_w3288_v;
	wire v_w1892_v;
	wire v_w4033_v;
	wire v_w5142_v;
	reg v_s347_v;
	wire v_w4381_v;
	wire v_w8185_v;
	wire v_w3160_v;
	wire v_w5745_v;
	wire v_w4633_v;
	wire v_w6860_v;
	reg v_s171_v;
	wire v_w2620_v;
	wire v_w1636_v;
	wire v_w6325_v;
	wire v_w6872_v;
	wire v_w7351_v;
	wire v_w4923_v;
	wire v_w8022_v;
	wire v_w2169_v;
	wire v_w3051_v;
	wire v_w6900_v;
	wire v_w3148_v;
	wire v_w4240_v;
	wire v_w3560_v;
	wire v_w160_v;
	wire v_w1063_v;
	reg v_s497_v;
	wire v_w1032_v;
	wire v_w2621_v;
	wire v_w5001_v;
	wire v_w2367_v;
	wire v_w6559_v;
	wire v_w2373_v;
	wire v_w6868_v;
	wire v_w5190_v;
	wire v_w4788_v;
	wire v_w2384_v;
	wire v_w6418_v;
	wire v_w6041_v;
	wire v_w2579_v;
	wire v_w3447_v;
	wire v_w214_v;
	wire v_w3131_v;
	wire v_w2220_v;
	wire v_w3490_v;
	wire v_w3095_v;
	reg v_s322_v;
	wire v_w5915_v;
	wire v_w764_v;
	wire v_w3327_v;
	wire v_w1150_v;
	wire v_w7863_v;
	wire v_w359_v;
	wire v_w3953_v;
	wire v_w4124_v;
	wire v_w4678_v;
	wire v_w6994_v;
	wire v_w3876_v;
	wire v_w5401_v;
	wire v_w3579_v;
	wire v_w2067_v;
	wire v_w7079_v;
	wire v_w1500_v;
	wire v_w4116_v;
	wire v_w2276_v;
	wire v_w6411_v;
	wire v_w2200_v;
	reg v_s372_v;
	wire v_w3820_v;
	wire v_w4997_v;
	reg v_s101_v;
	wire v_w6822_v;
	wire v_w6807_v;
	wire v_w7300_v;
	wire v_w2398_v;
	wire v_w3002_v;
	wire v_w3340_v;
	wire v_w99_v;
	wire v_w193_v;
	reg v_s155_v;
	wire v_w8212_v;
	reg v_s188_v;
	wire v_w6425_v;
	wire v_w1275_v;
	wire v_w1229_v;
	wire v_w780_v;
	wire v_w4676_v;
	wire v_w1169_v;
	wire v_w2250_v;
	wire v_w5623_v;
	wire v_w2634_v;
	wire v_w689_v;
	wire v_w3103_v;
	wire v_w1763_v;
	wire v_w7259_v;
	wire v_w5589_v;
	wire v_w6015_v;
	wire v_w7470_v;
	wire v_w4605_v;
	wire v_w194_v;
	wire v_w1945_v;
	wire v_w1538_v;
	wire v_w3763_v;
	wire v_w2914_v;
	wire v_w3753_v;
	wire v_w3887_v;
	wire v_w3502_v;
	wire v_w2858_v;
	wire v_w3918_v;
	wire v_w4439_v;
	wire v_w8060_v;
	wire v_w325_v;
	wire v_w7159_v;
	wire v_w4819_v;
	wire v_w259_v;
	wire v_w3875_v;
	wire v_w1124_v;
	wire v_w1776_v;
	wire v_w2627_v;
	wire v_w3496_v;
	wire v_w7340_v;
	wire v_w1761_v;
	wire v_w548_v;
	wire v_w6899_v;
	wire v_w1428_v;
	wire v_w5024_v;
	wire v_w604_v;
	wire v_w3232_v;
	reg v_s332_v;
	wire v_w5307_v;
	wire v_w4989_v;
	wire v_w1348_v;
	wire v_w6647_v;
	wire v_w2595_v;
	wire v_w4245_v;
	wire v_w2305_v;
	wire v_w6840_v;
	wire v_w1715_v;
	wire v_w483_v;
	wire v_w8108_v;
	wire v_w4201_v;
	wire v_w3799_v;
	wire v_w4413_v;
	wire v_w2438_v;
	wire v_w7453_v;
	wire v_w7970_v;
	wire v_w6499_v;
	wire v_w208_v;
	wire v_w5901_v;
	wire v_w4862_v;
	wire v_w3800_v;
	wire v_w1293_v;
	wire v_w602_v;
	reg v_s73_v;
	reg v_s148_v;
	wire v_w4102_v;
	wire v_w6328_v;
	wire v_w7668_v;
	wire v_w6769_v;
	wire v_w7742_v;
	wire v_w131_v;
	wire v_w4510_v;
	wire v_w7647_v;
	wire v_w8167_v;
	wire v_w7984_v;
	wire v_w5347_v;
	wire v_w5835_v;
	wire v_w6162_v;
	wire v_w4907_v;
	wire v_w2531_v;
	wire v_w6283_v;
	wire v_w7172_v;
	wire v_w5847_v;
	wire v_w5724_v;
	wire v_w5406_v;
	wire v_w3809_v;
	wire v_w424_v;
	reg v_s84_v;
	wire v_w1181_v;
	wire v_w2295_v;
	reg v_s469_v;
	wire v_w3383_v;
	wire v_w6606_v;
	wire v_w4990_v;
	reg v_s301_v;
	wire v_w352_v;
	wire v_w4312_v;
	wire v_w8075_v;
	wire v_w6392_v;
	reg v_s176_v;
	wire v_w2738_v;
	wire v_w3717_v;
	wire v_w486_v;
	wire v_w6_v;
	wire v_w6123_v;
	wire v_w6751_v;
	wire v_w5305_v;
	wire v_w4384_v;
	wire v_w4374_v;
	wire v_w4056_v;
	wire v_w5655_v;
	wire v_w989_v;
	wire v_w7382_v;
	wire v_w6029_v;
	wire v_w4755_v;
	wire v_w5702_v;
	wire v_w3601_v;
	wire v_w1376_v;
	wire v_w881_v;
	wire v_w2973_v;
	wire v_w7271_v;
	wire v_w5557_v;
	wire v_w390_v;
	wire v_w5168_v;
	wire v_w4254_v;
	wire v_w188_v;
	wire v_w3909_v;
	wire v_w879_v;
	wire v_w5193_v;
	wire v_w111_v;
	wire v_w1112_v;
	wire v_w6591_v;
	wire v_w4110_v;
	wire v_w733_v;
	wire v_w7661_v;
	wire v_w2722_v;
	wire v_w6024_v;
	reg v_s345_v;
	wire v_w2287_v;
	wire v_w4322_v;
	reg v_s58_v;
	wire v_w8100_v;
	wire v_w6168_v;
	wire v_w1278_v;
	wire v_w7956_v;
	wire v_w5108_v;
	wire v_w5794_v;
	wire v_w7030_v;
	reg v_s143_v;
	wire v_w7334_v;
	wire v_w657_v;
	wire v_w7697_v;
	wire v_w3903_v;
	wire v_w2687_v;
	wire v_w7601_v;
	wire v_w4596_v;
	wire v_w6703_v;
	wire v_w4921_v;
	wire v_w6657_v;
	wire v_w5948_v;
	wire v_w6747_v;
	wire v_w2834_v;
	wire v_w7337_v;
	wire v_w5464_v;
	wire v_w205_v;
	wire v_w143_v;
	wire v_w4095_v;
	wire v_w7423_v;
	wire v_w3834_v;
	wire v_w4951_v;
	reg v_s386_v;
	wire v_w7655_v;
	wire v_w7074_v;
	wire v_w5304_v;
	wire v_w7853_v;
	wire v_w5112_v;
	wire v_w7820_v;
	wire v_w6605_v;
	wire v_w2783_v;
	wire v_w117_v;
	wire v_w2588_v;
	wire v_w6616_v;
	wire v_w2793_v;
	wire v_w3668_v;
	wire v_w6167_v;
	wire v_w6092_v;
	wire v_w3557_v;
	wire v_w6595_v;
	wire v_w4062_v;
	wire v_w1355_v;
	reg v_s427_v;
	wire v_w1317_v;
	wire v_w4912_v;
	wire v_w7792_v;
	wire v_w3033_v;
	wire v_w6575_v;
	wire v_w942_v;
	wire v_w4537_v;
	wire v_w1328_v;
	reg v_s159_v;
	wire v_w6216_v;
	wire v_w2565_v;
	wire v_w2585_v;
	wire v_w4182_v;
	wire v_w438_v;
	wire v_w6478_v;
	wire v_w8073_v;
	wire v_w2159_v;
	wire v_w800_v;
	wire v_w2291_v;
	wire v_w1879_v;
	wire v_w6627_v;
	wire v_w6503_v;
	wire v_w912_v;
	reg v_s12_v;
	wire v_w7940_v;
	wire v_w306_v;
	wire v_w5620_v;
	wire v_w5048_v;
	wire v_w7176_v;
	wire v_w778_v;
	wire v_w815_v;
	wire v_w2658_v;
	wire v_w5996_v;
	wire v_w7451_v;
	wire v_w1579_v;
	wire v_w7452_v;
	wire v_w1811_v;
	wire v_w5629_v;
	wire v_w1969_v;
	wire v_w5549_v;
	wire v_w506_v;
	wire v_w3534_v;
	wire v_w3645_v;
	wire v_w10_v;
	wire v_w5405_v;
	wire v_w3781_v;
	wire v_w8036_v;
	reg v_s16_v;
	wire v_w417_v;
	wire v_w7481_v;
	wire v_w4277_v;
	wire v_w6734_v;
	wire v_w4144_v;
	wire v_w6848_v;
	wire v_w7004_v;
	wire v_w3863_v;
	wire v_w5720_v;
	wire v_w1557_v;
	wire v_w8015_v;
	wire v_w140_v;
	wire v_w2647_v;
	wire v_w3083_v;
	wire v_w2855_v;
	wire v_w7272_v;
	wire v_w5211_v;
	wire v_w1218_v;
	wire v_w5035_v;
	wire v_w5849_v;
	wire v_w3839_v;
	reg v_s74_v;
	wire v_w1924_v;
	wire v_w3529_v;
	wire v_w3760_v;
	wire v_w7732_v;
	wire v_w6871_v;
	wire v_w6794_v;
	wire v_w1437_v;
	wire v_w4043_v;
	wire v_w6897_v;
	reg v_s452_v;
	wire v_w1140_v;
	wire v_w1459_v;
	wire v_w596_v;
	wire v_w4942_v;
	wire v_w671_v;
	wire v_w4524_v;
	wire v_w1807_v;
	wire v_w3238_v;
	wire v_w5555_v;
	reg v_s460_v;
	wire v_w2781_v;
	wire v_w5505_v;
	wire v_w770_v;
	wire v_w4617_v;
	wire v_w4198_v;
	wire v_w4947_v;
	wire v_w6145_v;
	wire v_w4368_v;
	wire v_w7983_v;
	wire v_w4785_v;
	wire v_w4936_v;
	wire v_w5869_v;
	reg v_s37_v;
	wire v_w1062_v;
	wire v_w260_v;
	wire v_w5019_v;
	wire v_w968_v;
	wire v_w7352_v;
	wire v_w1382_v;
	wire v_w7842_v;
	wire v_w1188_v;
	wire v_w4434_v;
	wire v_w219_v;
	wire v_w8031_v;
	wire v_w832_v;
	wire v_w430_v;
	wire v_w2272_v;
	wire v_w6620_v;
	wire v_w1865_v;
	wire v_w4653_v;
	wire v_w1549_v;
	wire v_w2718_v;
	wire v_w2279_v;
	wire v_w4387_v;
	wire v_w2697_v;
	wire v_w712_v;
	wire v_w5658_v;
	wire v_w5742_v;
	wire v_w5554_v;
	wire v_w3906_v;
	wire v_w7433_v;
	wire v_w3929_v;
	wire v_w5562_v;
	wire v_w5467_v;
	wire v_w4825_v;
	wire v_w2418_v;
	wire v_w8156_v;
	wire v_w1116_v;
	reg v_s131_v;
	wire v_w6511_v;
	wire v_w7645_v;
	wire v_w385_v;
	wire v_w3582_v;
	wire v_w4337_v;
	wire v_w8027_v;
	wire v_w5319_v;
	wire v_w4539_v;
	wire v_w5744_v;
	wire v_w1192_v;
	reg v_s421_v;
	wire v_w7329_v;
	wire v_w6737_v;
	reg v_s233_v;
	wire v_w7579_v;
	wire v_w6379_v;
	wire v_w509_v;
	wire v_w5568_v;
	wire v_w2473_v;
	wire v_w6281_v;
	wire v_w1767_v;
	wire v_w1605_v;
	wire v_w5110_v;
	wire v_w1228_v;
	wire v_w4574_v;
	wire v_w6801_v;
	wire v_w1773_v;
	wire v_w6623_v;
	wire v_w5645_v;
	wire v_w5529_v;
	wire v_w5547_v;
	wire v_w1009_v;
	wire v_w3034_v;
	wire v_w6950_v;
	wire v_w723_v;
	wire v_w6208_v;
	reg v_s170_v;
	wire v_w5422_v;
	wire v_w754_v;
	wire v_w6587_v;
	wire v_w4843_v;
	wire v_w7869_v;
	wire v_w5771_v;
	wire v_w6484_v;
	wire v_w6684_v;
	wire v_w8038_v;
	wire v_w5992_v;
	wire v_w3305_v;
	wire v_w7495_v;
	wire v_w6829_v;
	wire v_w4999_v;
	wire v_w278_v;
	wire v_w4558_v;
	reg v_s162_v;
	wire v_w7435_v;
	wire v_w1626_v;
	wire v_w5264_v;
	wire v_w3249_v;
	wire v_w6686_v;
	wire v_w790_v;
	wire v_w2001_v;
	wire v_w7234_v;
	wire v_w3732_v;
	wire v_w395_v;
	wire v_w759_v;
	reg v_s416_v;
	wire v_w2592_v;
	wire v_w1677_v;
	wire v_w5084_v;
	wire v_w1864_v;
	reg v_s52_v;
	wire v_w4363_v;
	wire v_w1615_v;
	wire v_w2307_v;
	wire v_w4067_v;
	wire v_w2198_v;
	wire v_w7714_v;
	wire v_w701_v;
	wire v_w2360_v;
	wire v_w4150_v;
	wire v_w1252_v;
	wire v_w59_v;
	wire v_w5261_v;
	wire v_w7816_v;
	wire v_w2417_v;
	wire v_w2773_v;
	wire v_w866_v;
	wire v_w698_v;
	wire v_w6020_v;
	wire v_w3631_v;
	reg v_s33_v;
	wire v_w2230_v;
	reg v_s46_v;
	wire v_w3405_v;
	wire v_w4467_v;
	wire v_w2529_v;
	wire v_w7160_v;
	wire v_w7293_v;
	wire v_w5281_v;
	wire v_w4141_v;
	wire v_w3765_v;
	wire v_w2033_v;
	wire v_w8142_v;
	wire v_w4053_v;
	wire v_w150_v;
	wire v_w3217_v;
	wire v_w6563_v;
	wire v_w7199_v;
	wire v_w6758_v;
	wire v_w7022_v;
	wire v_w4461_v;
	wire v_w7849_v;
	reg v_s473_v;
	wire v_w1933_v;
	wire v_w2583_v;
	wire v_w1870_v;
	wire v_w16_v;
	wire v_w6446_v;
	wire v_w5700_v;
	wire v_w2525_v;
	wire v_w2678_v;
	wire v_w7422_v;
	wire v_w3030_v;
	wire v_w7036_v;
	wire v_w2429_v;
	wire v_w6743_v;
	wire v_w4321_v;
	wire v_w900_v;
	wire v_w6967_v;
	wire v_w1154_v;
	wire v_w7562_v;
	wire v_w738_v;
	wire v_w2251_v;
	wire v_w6196_v;
	wire v_w7170_v;
	wire v_w386_v;
	wire v_w1312_v;
	wire v_w680_v;
	reg v_s361_v;
	wire v_w674_v;
	wire v_w5210_v;
	wire v_w5090_v;
	wire v_w6884_v;
	wire v_w1858_v;
	wire v_w1611_v;
	wire v_w1937_v;
	wire v_w1203_v;
	wire v_w4480_v;
	wire v_w5445_v;
	wire v_w316_v;
	reg v_s319_v;
	wire v_w6481_v;
	wire v_w7131_v;
	wire v_w4651_v;
	reg v_s376_v;
	wire v_w4642_v;
	wire v_w2976_v;
	wire v_w7006_v;
	wire v_w1282_v;
	wire v_w619_v;
	wire v_w3870_v;
	wire v_w4487_v;
	wire v_w1712_v;
	wire v_w4879_v;
	wire v_w236_v;
	wire v_w2511_v;
	wire v_w289_v;
	wire v_w1208_v;
	reg v_s178_v;
	wire v_w6841_v;
	wire v_w4995_v;
	wire v_w5581_v;
	wire v_w7325_v;
	wire v_w1489_v;
	wire v_w4531_v;
	wire v_w6072_v;
	wire v_w6368_v;
	wire v_w637_v;
	wire v_w6809_v;
	wire v_w2445_v;
	wire v_w7194_v;
	wire v_w3602_v;
	wire v_w945_v;
	reg v_s317_v;
	wire v_w5638_v;
	wire v_w2343_v;
	wire v_w2694_v;
	wire v_w822_v;
	wire v_w3444_v;
	wire v_w4269_v;
	wire v_w6908_v;
	wire v_w7828_v;
	reg v_s300_v;
	wire v_w1525_v;
	wire v_w3442_v;
	wire v_w3551_v;
	reg v_s119_v;
	wire v_w6991_v;
	wire v_w4225_v;
	reg v_s75_v;
	wire v_w2241_v;
	wire v_w6546_v;
	wire v_w6393_v;
	wire v_w4905_v;
	wire v_w7274_v;
	wire v_w5164_v;
	wire v_w3312_v;
	wire v_w4013_v;
	wire v_w1418_v;
	wire v_w4650_v;
	wire v_w5100_v;
	wire v_w7232_v;
	wire v_w6704_v;
	wire v_w3818_v;
	wire v_w7333_v;
	wire v_w7248_v;
	wire v_w6593_v;
	wire v_w8078_v;
	wire v_w8218_v;
	wire v_w2441_v;
	wire v_w2638_v;
	wire v_w3628_v;
	wire v_w5689_v;
	wire v_w5293_v;
	reg v_s298_v;
	wire v_w6526_v;
	wire v_w1344_v;
	wire v_w1245_v;
	wire v_w6726_v;
	wire v_w4959_v;
	wire v_w6492_v;
	wire v_w3945_v;
	wire v_w4656_v;
	wire v_w760_v;
	wire v_w6125_v;
	wire v_w4697_v;
	wire v_w286_v;
	wire v_w3605_v;
	wire v_w7851_v;
	wire v_o18_v;
	wire v_w7494_v;
	wire v_w5071_v;
	wire v_w2171_v;
	wire v_w1744_v;
	wire v_w4313_v;
	wire v_w3248_v;
	wire v_w7787_v;
	wire v_w4154_v;
	wire v_w2102_v;
	wire v_w4283_v;
	wire v_w4304_v;
	wire v_w7929_v;
	wire v_w5971_v;
	wire v_w6570_v;
	wire v_w3074_v;
	wire v_w435_v;
	wire v_w2546_v;
	wire v_w1171_v;
	wire v_w7631_v;
	wire v_w2216_v;
	wire v_w7744_v;
	wire v_w1397_v;
	wire v_w4750_v;
	wire v_w4472_v;
	wire v_w6157_v;
	wire v_w3804_v;
	wire v_w2504_v;
	wire v_w3563_v;
	wire v_w7357_v;
	wire v_w2165_v;
	wire v_w1274_v;
	wire v_w5808_v;
	reg v_s373_v;
	wire v_w7123_v;
	wire v_w4089_v;
	wire v_w4230_v;
	wire v_w3419_v;
	wire v_w4042_v;
	wire v_w4762_v;
	wire v_w632_v;
	reg v_s401_v;
	wire v_w5141_v;
	wire v_w135_v;
	wire v_w3158_v;
	wire v_w5105_v;
	wire v_w5381_v;
	wire v_w1132_v;
	wire v_w1859_v;
	wire v_w7882_v;
	wire v_w5768_v;
	wire v_w7814_v;
	reg v_s480_v;
	wire v_w6655_v;
	wire v_w5600_v;
	wire v_w6428_v;
	wire v_w1241_v;
	wire v_w18_v;
	wire v_w5811_v;
	wire v_w1223_v;
	wire v_w6700_v;
	wire v_w6488_v;
	wire v_w2505_v;
	wire v_w3741_v;
	wire v_w7258_v;
	wire v_w4227_v;
	wire v_w239_v;
	wire v_w2887_v;
	wire v_w5286_v;
	wire v_w243_v;
	wire v_w995_v;
	reg v_s234_v;
	wire v_w661_v;
	wire v_w3063_v;
	wire v_w3568_v;
	wire v_w890_v;
	wire v_w8057_v;
	wire v_w5348_v;
	wire v_w6226_v;
	wire v_w4106_v;
	wire v_w6271_v;
	wire v_w6919_v;
	wire v_w1139_v;
	wire v_w1238_v;
	wire v_w387_v;
	wire v_w7810_v;
	wire v_w5393_v;
	wire v_w3743_v;
	wire v_w8063_v;
	wire v_w473_v;
	wire v_w576_v;
	wire v_w6084_v;
	wire v_w6455_v;
	wire v_w757_v;
	wire v_w7067_v;
	wire v_w3736_v;
	wire v_w2232_v;
	wire v_w5649_v;
	wire v_w420_v;
	wire v_w1556_v;
	wire v_w5591_v;
	wire v_w2231_v;
	wire v_w109_v;
	wire v_w2829_v;
	wire v_w978_v;
	wire v_w304_v;
	wire v_w5934_v;
	wire v_w5532_v;
	wire v_w2106_v;
	wire v_w591_v;
	wire v_w818_v;
	reg v_s135_v;
	wire v_w4064_v;
	reg v_s41_v;
	wire v_w5598_v;
	wire v_w1237_v;
	wire v_w1294_v;
	wire v_w2166_v;
	wire v_w4267_v;
	wire v_w813_v;
	wire v_w5397_v;
	wire v_w5427_v;
	wire v_w2557_v;
	wire v_w5385_v;
	wire v_w6381_v;
	wire v_w1804_v;
	wire v_w739_v;
	wire v_w2882_v;
	wire v_w4133_v;
	wire v_w4405_v;
	wire v_w4169_v;
	wire v_w4291_v;
	wire v_w3704_v;
	wire v_w481_v;
	wire v_w4584_v;
	wire v_w3626_v;
	wire v_w5991_v;
	wire v_w7307_v;
	wire v_w4647_v;
	wire v_w4764_v;
	wire v_w53_v;
	wire v_w4877_v;
	wire v_w7871_v;
	wire v_w7317_v;
	wire v_w7745_v;
	wire v_w7884_v;
	wire v_w5718_v;
	wire v_w4552_v;
	wire v_w3984_v;
	wire v_w130_v;
	wire v_w1654_v;
	wire v_w1349_v;
	wire v_w455_v;
	wire v_w7663_v;
	wire v_w1943_v;
	wire v_w6996_v;
	wire v_w1652_v;
	wire v_w170_v;
	wire v_w5236_v;
	wire v_w6589_v;
	wire v_w8244_v;
	wire v_w1054_v;
	wire v_w835_v;
	wire v_w5756_v;
	wire v_w4433_v;
	wire v_w7941_v;
	wire v_w7746_v;
	wire v_w777_v;
	wire v_w153_v;
	wire v_w3292_v;
	wire v_w5905_v;
	wire v_w4556_v;
	wire v_w3853_v;
	wire v_w3070_v;
	wire v_w6586_v;
	wire v_w3888_v;
	wire v_w1195_v;
	wire v_w4176_v;
	wire v_w4449_v;
	wire v_w4037_v;
	wire v_w1760_v;
	wire v_w7684_v;
	wire v_w1010_v;
	wire v_w296_v;
	wire v_w4661_v;
	wire v_w2432_v;
	wire v_w8182_v;
	wire v_w6752_v;
	wire v_w3932_v;
	wire v_w5959_v;
	wire v_w5545_v;
	wire v_w3380_v;
	wire v_w5075_v;
	reg v_s260_v;
	reg v_s430_v;
	wire v_w6881_v;
	wire v_w1077_v;
	wire v_w4465_v;
	wire v_w5109_v;
	wire v_w4162_v;
	wire v_w5714_v;
	wire v_w2375_v;
	wire v_w4323_v;
	wire v_w915_v;
	wire v_w2806_v;
	wire v_w1918_v;
	wire v_w5136_v;
	wire v_w1176_v;
	wire v_w1134_v;
	wire v_w6865_v;
	wire v_w1794_v;
	wire v_w3613_v;
	wire v_w7753_v;
	wire v_w725_v;
	reg v_s329_v;
	wire v_w1868_v;
	wire v_w2013_v;
	wire v_w4431_v;
	wire v_w2630_v;
	wire v_w1766_v;
	reg v_s134_v;
	wire v_w1287_v;
	wire v_w5368_v;
	wire v_w1915_v;
	wire v_w500_v;
	wire v_w6335_v;
	wire v_w5080_v;
	wire v_w6641_v;
	wire v_w1213_v;
	wire v_w4735_v;
	wire v_w5778_v;
	wire v_w2597_v;
	wire v_w1873_v;
	wire v_w298_v;
	wire v_w1703_v;
	wire v_w834_v;
	wire v_w7260_v;
	wire v_w552_v;
	wire v_w3565_v;
	wire v_w4021_v;
	reg v_s350_v;
	wire v_w327_v;
	wire v_w2852_v;
	wire v_w6456_v;
	wire v_w662_v;
	wire v_w4356_v;
	wire v_w4071_v;
	wire v_w6750_v;
	wire v_w2093_v;
	wire v_w1511_v;
	wire v_w4545_v;
	wire v_w7449_v;
	wire v_w8195_v;
	wire v_w23_v;
	wire v_w6242_v;
	wire v_w639_v;
	wire v_w3307_v;
	wire v_w819_v;
	wire v_w141_v;
	wire v_w2470_v;
	wire v_w1120_v;
	wire v_w2321_v;
	wire v_w1501_v;
	wire v_w5499_v;
	wire v_w2843_v;
	reg v_s202_v;
	wire v_w4305_v;
	wire v_w3381_v;
	wire v_w4813_v;
	reg v_s50_v;
	wire v_w1304_v;
	wire v_w7011_v;
	wire v_w1184_v;
	wire v_w1297_v;
	wire v_w3049_v;
	wire v_w1187_v;
	wire v_w5796_v;
	wire v_w464_v;
	wire v_w7501_v;
	wire v_w469_v;
	wire v_w3538_v;
	wire v_w8093_v;
	wire v_w3493_v;
	wire v_w5608_v;
	wire v_w1224_v;
	wire v_w1512_v;
	wire v_w7829_v;
	wire v_w1488_v;
	wire v_w847_v;
	wire v_w3756_v;
	wire v_w1625_v;
	wire v_w7972_v;
	wire v_w2076_v;
	wire v_w6744_v;
	wire v_w7767_v;
	wire v_w6768_v;
	wire v_w4566_v;
	wire v_w1455_v;
	wire v_w1507_v;
	wire v_w3263_v;
	wire v_w4823_v;
	wire v_w2126_v;
	wire v_w3997_v;
	wire v_w4731_v;
	wire v_w5188_v;
	reg v_s181_v;
	wire v_w6934_v;
	wire v_w3933_v;
	wire v_w4627_v;
	reg v_s316_v;
	wire v_w946_v;
	wire v_w282_v;
	wire v_w7537_v;
	wire v_w2667_v;
	wire v_w926_v;
	wire v_w4869_v;
	wire v_w635_v;
	wire v_w3151_v;
	wire v_w7332_v;
	wire v_w3609_v;
	reg v_s338_v;
	wire v_w934_v;
	reg v_s501_v;
	wire v_w3793_v;
	wire v_w6678_v;
	wire v_w2791_v;
	wire v_w6032_v;
	wire v_w1029_v;
	reg v_s220_v;
	wire v_w7064_v;
	wire v_w735_v;
	wire v_w3367_v;
	wire v_w4324_v;
	wire v_w6864_v;
	wire v_w8190_v;
	wire v_w3455_v;
	wire v_w4564_v;
	reg v_s201_v;
	wire v_w3691_v;
	wire v_w5309_v;
	wire v_w2333_v;
	wire v_w3780_v;
	wire v_w5734_v;
	wire v_w2131_v;
	wire v_w7864_v;
	wire v_w2578_v;
	reg v_s315_v;
	wire v_w534_v;
	reg v_s243_v;
	wire v_w4931_v;
	wire v_w27_v;
	wire v_w419_v;
	wire v_w7936_v;
	wire v_w2709_v;
	wire v_w6982_v;
	wire v_w883_v;
	wire v_w2507_v;
	wire v_w2188_v;
	wire v_w1125_v;
	reg v_s125_v;
	wire v_w5686_v;
	wire v_w5040_v;
	wire v_w6134_v;
	reg v_s15_v;
	wire v_w2129_v;
	wire v_w2528_v;
	wire v_w2548_v;
	wire v_w5631_v;
	wire v_w7492_v;
	wire v_w5947_v;
	wire v_w6192_v;
	wire v_w830_v;
	wire v_w2935_v;
	wire v_w2696_v;
	wire v_w4974_v;
	wire v_w758_v;
	wire v_w39_v;
	wire v_w8126_v;
	wire v_w4723_v;
	wire v_w3971_v;
	wire v_w7890_v;
	wire v_w4380_v;
	wire v_w958_v;
	wire v_w782_v;
	wire v_w7759_v;
	wire v_w7775_v;
	wire v_w3318_v;
	wire v_w5824_v;
	wire v_w3420_v;
	wire v_w3202_v;
	reg v_s450_v;
	wire v_w4649_v;
	wire v_w5351_v;
	wire v_w7996_v;
	wire v_w2841_v;
	wire v_w2705_v;
	wire v_w1426_v;
	wire v_w3730_v;
	wire v_w1109_v;
	wire v_w1221_v;
	wire v_w5404_v;
	wire v_w6483_v;
	wire v_w1576_v;
	reg v_s310_v;
	wire v_w4576_v;
	wire v_w3738_v;
	wire v_w4076_v;
	wire v_w1903_v;
	reg v_s21_v;
	wire v_w5421_v;
	wire v_w1225_v;
	wire v_w5970_v;
	wire v_w4732_v;
	wire v_w954_v;
	wire v_w562_v;
	wire v_w6188_v;
	wire v_w7809_v;
	wire v_w7014_v;
	wire v_w5419_v;
	wire v_w4833_v;
	wire v_w1204_v;
	wire v_w4083_v;
	wire v_w7255_v;
	wire v_w5922_v;
	wire v_w1709_v;
	wire v_w1276_v;
	wire v_w6399_v;
	wire v_w8089_v;
	wire v_w4643_v;
	wire v_w7187_v;
	wire v_w26_v;
	wire v_w7613_v;
	wire v_w1194_v;
	wire v_w3193_v;
	wire v_w2831_v;
	wire v_w5983_v;
	wire v_w5748_v;
	wire v_w1970_v;
	wire v_w6764_v;
	wire v_w2862_v;
	wire v_w5342_v;
	wire v_w7309_v;
	wire v_w6417_v;
	wire v_w5224_v;
	wire v_w7522_v;
	wire v_w5727_v;
	wire v_w2972_v;
	wire v_w6334_v;
	reg v_s76_v;
	wire v_w5617_v;
	wire v_w7902_v;
	wire v_w7376_v;
	wire v_w3513_v;
	wire v_w6332_v;
	wire v_w4000_v;
	wire v_w5708_v;
	wire v_w5833_v;
	wire v_w6293_v;
	wire v_w6317_v;
	wire v_w91_v;
	wire v_w3608_v;
	wire v_w4421_v;
	wire v_w3546_v;
	wire v_w7818_v;
	reg v_s311_v;
	wire v_w6185_v;
	wire v_w652_v;
	wire v_w6514_v;
	wire v_w1244_v;
	wire v_w3355_v;
	reg v_s357_v;
	wire v_w6378_v;
	wire v_w1100_v;
	wire v_w6540_v;
	wire v_w4253_v;
	wire v_w6078_v;
	wire v_w7412_v;
	wire v_w801_v;
	wire v_w6479_v;
	wire v_w2629_v;
	wire v_w6988_v;
	wire v_w4127_v;
	wire v_w6272_v;
	wire v_w2784_v;
	reg v_s463_v;
	wire v_w5396_v;
	wire v_w1291_v;
	wire v_w1745_v;
	wire v_w542_v;
	wire v_w5266_v;
	wire v_w5115_v;
	wire v_w2981_v;
	wire v_w3372_v;
	wire v_w4035_v;
	wire v_w5885_v;
	wire v_w4496_v;
	wire v_w785_v;
	wire v_w8018_v;
	wire v_w1529_v;
	wire v_w8191_v;
	wire v_w3413_v;
	wire v_w4122_v;
	wire v_w3366_v;
	wire v_w3890_v;
	wire v_w1069_v;
	wire v_w4244_v;
	wire v_w7402_v;
	wire v_w3564_v;
	wire v_w4261_v;
	wire v_w4726_v;
	wire v_w2666_v;
	wire v_w1629_v;
	wire v_w4855_v;
	wire v_w3394_v;
	wire v_w5647_v;
	wire v_w6772_v;
	wire v_w3235_v;
	wire v_w2488_v;
	reg v_s312_v;
	wire v_w1391_v;
	wire v_w1453_v;
	wire v_w2735_v;
	wire v_w3951_v;
	wire v_w1881_v;
	wire v_w6438_v;
	wire v_w4847_v;
	wire v_w1085_v;
	wire v_w6388_v;
	wire v_w979_v;
	wire v_w2246_v;
	wire v_w6326_v;
	wire v_w5098_v;
	wire v_w1505_v;
	wire v_w7538_v;
	wire v_w443_v;
	wire v_w1648_v;
	wire v_w183_v;
	wire v_w590_v;
	wire v_w7285_v;
	wire v_w7049_v;
	wire v_w3878_v;
	wire v_w6444_v;
	wire v_w5508_v;
	wire v_w728_v;
	wire v_w3777_v;
	wire v_w6221_v;
	wire v_w544_v;
	wire v_w361_v;
	wire v_w4178_v;
	wire v_w2335_v;
	wire v_w3549_v;
	wire v_w2856_v;
	wire v_w5237_v;
	wire v_w4828_v;
	wire v_w1706_v;
	wire v_w8227_v;
	wire v_w4674_v;
	wire v_w8254_v;
	wire v_w7901_v;
	wire v_w5838_v;
	wire v_w4077_v;
	wire v_w1086_v;
	reg v_s360_v;
	wire v_w6630_v;
	wire v_w4771_v;
	wire v_w3595_v;
	wire v_w2746_v;
	wire v_w8072_v;
	wire v_w8023_v;
	wire v_w6666_v;
	wire v_w5219_v;
	wire v_w539_v;
	wire v_w831_v;
	wire v_w6111_v;
	wire v_w616_v;
	wire v_w7948_v;
	reg v_s465_v;
	wire v_w4512_v;
	wire v_w6594_v;
	wire v_w3745_v;
	wire v_w5063_v;
	wire v_w1156_v;
	wire v_w3998_v;
	wire v_w7386_v;
	wire v_w3254_v;
	wire v_w1445_v;
	wire v_w2676_v;
	wire v_w7727_v;
	wire v_w7429_v;
	wire v_w4262_v;
	wire v_w948_v;
	wire v_w7805_v;
	wire v_w440_v;
	wire v_w4822_v;
	wire v_w8008_v;
	wire v_w5584_v;
	wire v_w5488_v;
	wire v_w1060_v;
	wire v_w334_v;
	wire v_w3517_v;
	wire v_w6879_v;
	wire v_w5531_v;
	wire v_w6096_v;
	wire v_w1309_v;
	wire v_w3007_v;
	wire v_w4725_v;
	wire v_w2698_v;
	wire v_w1535_v;
	wire v_w2601_v;
	wire v_w8209_v;
	wire v_w7958_v;
	wire v_w3621_v;
	wire v_w5214_v;
	reg v_s381_v;
	wire v_w457_v;
	wire v_w5324_v;
	wire v_w1578_v;
	wire v_w80_v;
	wire v_w7565_v;
	wire v_w6017_v;
	wire v_w5717_v;
	wire v_w4386_v;
	wire v_w4543_v;
	wire v_w1185_v;
	wire v_w7604_v;
	wire v_w4623_v;
	wire v_w300_v;
	wire v_w5988_v;
	wire v_w2616_v;
	wire v_w4286_v;
	wire v_w6846_v;
	wire v_w6845_v;
	wire v_w5262_v;
	wire v_w1353_v;
	wire v_w6981_v;
	wire v_w3501_v;
	wire v_w7935_v;
	wire v_w6007_v;
	wire v_w3416_v;
	wire v_w3824_v;
	wire v_w5101_v;
	wire v_w7321_v;
	wire v_w6624_v;
	wire v_w4483_v;
	wire v_w4860_v;
	wire v_w574_v;
	wire v_w1388_v;
	wire v_w2758_v;
	wire v_w6174_v;
	wire v_w3308_v;
	wire v_w7254_v;
	wire v_w6918_v;
	wire v_w554_v;
	wire v_w851_v;
	wire v_w32_v;
	wire v_w5834_v;
	reg v_s224_v;
	wire v_w2741_v;
	wire v_w5990_v;
	wire v_w6956_v;
	wire v_w1517_v;
	wire v_w6873_v;
	wire v_w917_v;
	wire v_w2107_v;
	wire v_w6548_v;
	wire v_w70_v;
	wire v_w2606_v;
	wire v_w3640_v;
	wire v_w5276_v;
	wire v_w3230_v;
	wire v_w2364_v;
	wire v_w3247_v;
	wire v_w1680_v;
	wire v_w2436_v;
	wire v_w362_v;
	reg v_s391_v;
	reg v_s519_v;
	wire v_w4919_v;
	wire v_w4631_v;
	wire v_w5946_v;
	wire v_w7709_v;
	wire v_w3337_v;
	wire v_w423_v;
	wire v_w1016_v;
	wire v_w3556_v;
	wire v_w6672_v;
	wire v_w1262_v;
	wire v_w679_v;
	wire v_w4677_v;
	wire v_w1682_v;
	wire v_w4126_v;
	wire v_w3764_v;
	wire v_w2602_v;
	wire v_w8144_v;
	wire v_w4920_v;
	wire v_w157_v;
	wire v_w7676_v;
	wire v_w1775_v;
	wire v_w6792_v;
	wire v_w3710_v;
	wire v_w2314_v;
	wire v_w1663_v;
	wire v_w6914_v;
	reg v_s110_v;
	wire v_w891_v;
	wire v_w5739_v;
	wire v_w4794_v;
	wire v_w4263_v;
	wire v_w5764_v;
	wire v_w4008_v;
	wire v_w7195_v;
	wire v_w2728_v;
	wire v_w1250_v;
	wire v_w5612_v;
	wire v_w261_v;
	wire v_w5802_v;
	wire v_w3816_v;
	wire v_w1395_v;
	wire v_w4808_v;
	wire v_w2584_v;
	wire v_w4622_v;
	wire v_w1338_v;
	reg v_s425_v;
	wire v_w1743_v;
	wire v_w2282_v;
	wire v_w5476_v;
	wire v_w5274_v;
	wire v_w7513_v;
	wire v_w5721_v;
	wire v_w2422_v;
	wire v_w4916_v;
	wire v_w6331_v;
	wire v_w3651_v;
	wire v_w1843_v;
	wire v_w4477_v;
	wire v_w1255_v;
	wire v_w8077_v;
	wire v_w4977_v;
	wire v_w4469_v;
	reg v_s239_v;
	wire v_w3398_v;
	wire v_w6861_v;
	wire v_w7200_v;
	wire v_w206_v;
	wire v_w1860_v;
	wire v_w2304_v;
	wire v_w3572_v;
	wire v_w6902_v;
	reg v_s441_v;
	reg v_s333_v;
	wire v_w4657_v;
	wire v_w1479_v;
	wire v_w3889_v;
	wire v_w3452_v;
	wire v_w6898_v;
	wire v_w844_v;
	wire v_w1959_v;
	wire v_w6611_v;
	wire v_w2055_v;
	wire v_w3241_v;
	wire v_w624_v;
	wire v_w4460_v;
	wire v_w4355_v;
	wire v_w7974_v;
	wire v_w5513_v;
	wire v_w2506_v;
	wire v_w2493_v;
	wire v_w6246_v;
	wire v_w2091_v;
	wire v_w7789_v;
	wire v_w3826_v;
	reg v_s1_v;
	wire v_w753_v;
	wire v_w7951_v;
	wire v_w235_v;
	wire v_w1155_v;
	wire v_w4885_v;
	wire v_w6948_v;
	wire v_w3771_v;
	wire v_w2815_v;
	wire v_w5359_v;
	wire v_w6896_v;
	wire v_w8245_v;
	wire v_w5183_v;
	wire v_w4851_v;
	wire v_w4969_v;
	wire v_w2757_v;
	wire v_w3526_v;
	wire v_w7462_v;
	wire v_w2448_v;
	wire v_w5863_v;
	wire v_w8041_v;
	wire v_w6513_v;
	wire v_w7997_v;
	wire v_w1104_v;
	wire v_w113_v;
	wire v_w693_v;
	wire v_w7060_v;
	wire v_w1411_v;
	wire v_w7705_v;
	wire v_w7207_v;
	wire v_w575_v;
	wire v_o13_v;
	wire v_w3550_v;
	wire v_w174_v;
	wire v_w4728_v;
	wire v_w33_v;
	wire v_w3453_v;
	wire v_w1474_v;
	reg v_s453_v;
	wire v_w6716_v;
	wire v_w3168_v;
	wire v_w5622_v;
	wire v_w3854_v;
	wire v_w1753_v;
	wire v_w2509_v;
	wire v_w6160_v;
	wire v_w5976_v;
	wire v_w4616_v;
	wire v_w7344_v;
	wire v_w6314_v;
	wire v_w5697_v;
	wire v_w8102_v;
	reg v_s335_v;
	wire v_w1497_v;
	wire v_w7575_v;
	wire v_w1620_v;
	reg v_s57_v;
	wire v_w7437_v;
	wire v_w2368_v;
	wire v_w3940_v;
	wire v_w7044_v;
	reg v_s200_v;
	wire v_w5334_v;
	wire v_w6496_v;
	wire v_w7390_v;
	wire v_w1408_v;
	wire v_w2826_v;
	wire v_w6009_v;
	wire v_w3910_v;
	wire v_w4383_v;
	wire v_w766_v;
	wire v_w5674_v;
	wire v_w291_v;
	wire v_w2051_v;
	wire v_w4193_v;
	wire v_w1985_v;
	wire v_w5602_v;
	wire v_w2570_v;
	wire v_w6069_v;
	wire v_w6423_v;
	wire v_w4665_v;
	wire v_w1364_v;
	wire v_w350_v;
	wire v_w207_v;
	wire v_w2462_v;
	wire v_w5792_v;
	wire v_w6714_v;
	wire v_w1021_v;
	reg v_s180_v;
	wire v_w6638_v;
	wire v_w4290_v;
	wire v_w1424_v;
	wire v_w877_v;
	wire v_w180_v;
	wire v_w5884_v;
	wire v_w379_v;
	wire v_w4016_v;
	wire v_w1550_v;
	wire v_w2708_v;
	wire v_w2523_v;
	wire v_w1836_v;
	wire v_w7845_v;
	wire v_w5837_v;
	wire v_w54_v;
	wire v_w6825_v;
	wire v_w45_v;
	wire v_w7418_v;
	wire v_w2277_v;
	wire v_w6268_v;
	wire v_w4515_v;
	wire v_w1827_v;
	reg v_s185_v;
	wire v_w1366_v;
	wire v_w220_v;
	wire v_w2284_v;
	wire v_w1015_v;
	wire v_w7208_v;
	wire v_w7971_v;
	reg v_s506_v;
	wire v_w5234_v;
	wire v_w6779_v;
	wire v_w4807_v;
	wire v_w5540_v;
	wire v_w3392_v;
	wire v_w2905_v;
	wire v_w7076_v;
	wire v_w902_v;
	wire v_w6040_v;
	wire v_w3062_v;
	reg v_s268_v;
	wire v_w3020_v;
	wire v_w1565_v;
	wire v_w1942_v;
	wire v_w3724_v;
	wire v_w1577_v;
	wire v_w688_v;
	wire v_w4800_v;
	wire v_w2034_v;
	wire v_w899_v;
	wire v_w179_v;
	wire v_w1848_v;
	wire v_w2853_v;
	wire v_w3884_v;
	wire v_w6387_v;
	wire v_w3968_v;
	wire v_w6464_v;
	wire v_w7598_v;
	wire v_w4334_v;
	wire v_w6583_v;
	wire v_w5278_v;
	reg v_s172_v;
	wire v_w5634_v;
	wire v_w4535_v;
	wire v_w467_v;
	wire v_w5667_v;
	wire v_w7363_v;
	wire v_w5664_v;
	wire v_w213_v;
	wire v_w5953_v;
	wire v_w7409_v;
	wire v_w4369_v;
	wire v_w2184_v;
	wire v_w7881_v;
	wire v_w8052_v;
	wire v_w7824_v;
	wire v_w5036_v;
	wire v_w3173_v;
	wire v_w6172_v;
	wire v_w3014_v;
	wire v_w678_v;
	wire v_w5221_v;
	wire v_w7587_v;
	wire v_w1289_v;
	wire v_w6613_v;
	wire v_w6275_v;
	wire v_w7338_v;
	wire v_w3373_v;
	wire v_w4927_v;
	wire v_w3999_v;
	wire v_w2786_v;
	wire v_w3831_v;
	wire v_w378_v;
	wire v_w2377_v;
	wire v_w5517_v;
	wire v_w1008_v;
	reg v_s70_v;
	wire v_w5975_v;
	wire v_w2814_v;
	wire v_w3627_v;
	wire v_w4497_v;
	wire v_w2680_v;
	reg v_s66_v;
	wire v_w2986_v;
	reg v_s502_v;
	wire v_w6965_v;
	wire v_w1768_v;
	wire v_w763_v;
	wire v_w1732_v;
	wire v_w2140_v;
	wire v_w5719_v;
	wire v_w5472_v;
	wire v_w275_v;
	wire v_w6065_v;
	wire v_w5364_v;
	wire v_w4839_v;
	wire v_w6788_v;
	wire v_o16_v;
	wire v_w4086_v;
	wire v_w4917_v;
	wire v_w2691_v;
	wire v_w1669_v;
	wire v_w4475_v;
	wire v_w6402_v;
	wire v_w1197_v;
	wire v_w3432_v;
	wire v_w2382_v;
	wire v_w1955_v;
	wire v_w4758_v;
	wire v_w4404_v;
	reg v_s284_v;
	wire v_w5139_v;
	wire v_w7713_v;
	wire v_w3892_v;
	wire v_w3655_v;
	wire v_w1441_v;
	wire v_w3819_v;
	wire v_w3897_v;
	wire v_w4523_v;
	wire v_w1563_v;
	wire v_w4589_v;
	wire v_w4522_v;
	wire v_w4063_v;
	wire v_w2639_v;
	wire v_w5747_v;
	wire v_w6952_v;
	wire v_w5073_v;
	wire v_w5656_v;
	wire v_w4559_v;
	wire v_w4705_v;
	wire v_w7942_v;
	wire v_w317_v;
	wire v_w6625_v;
	wire v_w1067_v;
	wire v_w1708_v;
	wire v_w7364_v;
	reg v_s228_v;
	wire v_w1439_v;
	wire v_w1944_v;
	wire v_w5875_v;
	wire v_w6469_v;
	wire v_w7387_v;
	wire v_w2614_v;
	wire v_w292_v;
	wire v_w1842_v;
	wire v_w1266_v;
	wire v_w1271_v;
	wire v_w403_v;
	wire v_w5705_v;
	wire v_w4341_v;
	wire v_w3696_v;
	wire v_w2369_v;
	reg v_s422_v;
	wire v_w7648_v;
	wire v_w1961_v;
	wire v_w7542_v;
	reg v_s303_v;
	wire v_w4824_v;
	wire v_w5157_v;
	wire v_w4901_v;
	wire v_w2727_v;
	wire v_w6681_v;
	wire v_w472_v;
	wire v_w6863_v;
	wire v_w2020_v;
	wire v_w40_v;
	wire v_w5881_v;
	wire v_w1573_v;
	wire v_w545_v;
	wire v_w13_v;
	wire v_w2366_v;
	reg v_s3_v;
	wire v_w841_v;
	wire v_w4372_v;
	wire v_w1452_v;
	wire v_w5641_v;
	wire v_w907_v;
	wire v_w5923_v;
	wire v_w6463_v;
	wire v_w3396_v;
	wire v_w3757_v;
	wire v_w6236_v;
	wire v_w6095_v;
	wire v_w4217_v;
	wire v_w1339_v;
	wire v_w3844_v;
	reg v_s328_v;
	wire v_w5417_v;
	wire v_w3729_v;
	wire v_w4147_v;
	wire v_w4196_v;
	wire v_w2535_v;
	wire v_w5683_v;
	wire v_w8247_v;
	wire v_w5897_v;
	wire v_w7233_v;
	wire v_w2300_v;
	reg v_s174_v;
	wire v_w181_v;
	wire v_w2950_v;
	wire v_w6296_v;
	wire v_w852_v;
	wire v_w4527_v;
	wire v_w4586_v;
	reg v_s225_v;
	wire v_w1396_v;
	wire v_w846_v;
	wire v_w1429_v;
	wire v_w996_v;
	reg v_s493_v;
	wire v_w4444_v;
	wire v_w2745_v;
	wire v_w7350_v;
	wire v_w7722_v;
	wire v_w5780_v;
	wire v_w4926_v;
	wire v_w3927_v;
	wire v_w1850_v;
	wire v_w3508_v;
	wire v_w3713_v;
	wire v_w4403_v;
	wire v_w3618_v;
	wire v_w5848_v;
	wire v_w6777_v;
	wire v_w5941_v;
	wire v_w6960_v;
	wire v_w5855_v;
	wire v_w3949_v;
	wire v_w1270_v;
	wire v_w6882_v;
	wire v_w4471_v;
	wire v_w5310_v;
	wire v_w3136_v;
	wire v_w2700_v;
	wire v_w3071_v;
	wire v_w4113_v;
	wire v_w7960_v;
	wire v_w8096_v;
	wire v_w8070_v;
	wire v_w1456_v;
	wire v_w6955_v;
	wire v_w3446_v;
	wire v_w8235_v;
	wire v_w6549_v;
	wire v_w4389_v;
	wire v_w5066_v;
	wire v_w3064_v;
	wire v_w3905_v;
	wire v_w4085_v;
	wire v_w6651_v;
	wire v_w559_v;
	wire v_w6762_v;
	reg v_s218_v;
	wire v_w6303_v;
	wire v_w3441_v;
	wire v_w2407_v;
	wire v_w4209_v;
	wire v_w5189_v;
	wire v_w4131_v;
	wire v_w4121_v;
	wire v_w3919_v;
	wire v_w1115_v;
	wire v_w7168_v;
	wire v_w5202_v;
	wire v_w3857_v;
	wire v_w1667_v;
	wire v_w4123_v;
	wire v_w949_v;
	wire v_w7769_v;
	wire v_w3581_v;
	wire v_w5058_v;
	wire v_w6477_v;
	reg v_s321_v;
	wire v_w2956_v;
	wire v_w7728_v;
	wire v_w2132_v;
	wire v_w7302_v;
	wire v_w7448_v;
	wire v_w1995_v;
	wire v_w795_v;
	wire v_w1574_v;
	wire v_w1292_v;
	wire v_w7802_v;
	wire v_w1762_v;
	wire v_w6165_v;
	wire v_w3376_v;
	wire v_w5336_v;
	wire v_w1447_v;
	wire v_w7715_v;
	reg v_s133_v;
	wire v_w1313_v;
	wire v_w7257_v;
	wire v_w5593_v;
	wire v_w5377_v;
	wire v_w6545_v;
	wire v_w7371_v;
	wire v_w1404_v;
	wire v_w2918_v;
	wire v_w647_v;
	wire v_w3659_v;
	wire v_w838_v;
	wire v_w3375_v;
	wire v_w5325_v;
	wire v_w7380_v;
	wire v_w1350_v;
	wire v_w2199_v;
	wire v_w4883_v;
	wire v_w2109_v;
	wire v_w5500_v;
	wire v_w3143_v;
	wire v_w4107_v;
	wire v_w8137_v;
	wire v_w3611_v;
	wire v_w5954_v;
	wire v_w6004_v;
	wire v_w6421_v;
	wire v_w6554_v;
	wire v_w776_v;
	wire v_w3993_v;
	wire v_w7893_v;
	wire v_w3599_v;
	wire v_w4005_v;
	wire v_w4423_v;
	wire v_w2713_v;
	wire v_w2663_v;
	wire v_w8231_v;
	wire v_w5006_v;
	wire v_w1341_v;
	wire v_w7567_v;
	wire v_w5770_v;
	wire v_w4326_v;
	wire v_w5822_v;
	wire v_w1420_v;
	wire v_w5977_v;
	wire v_w5551_v;
	wire v_w3102_v;
	wire v_w7476_v;
	reg v_s459_v;
	wire v_w3693_v;
	wire v_w1782_v;
	wire v_w747_v;
	wire v_w3986_v;
	wire v_w6209_v;
	wire v_w2153_v;
	wire v_w2142_v;
	wire v_w1659_v;
	wire v_w8216_v;
	wire v_w120_v;
	wire v_w5124_v;
	wire v_w7897_v;
	wire v_w525_v;
	reg v_s20_v;
	wire v_w5496_v;
	wire v_w901_v;
	wire v_w4373_v;
	wire v_w5637_v;
	wire v_w5133_v;
	wire v_w6190_v;
	wire v_w2536_v;
	reg v_s384_v;
	wire v_w7640_v;
	wire v_w6181_v;
	wire v_w4853_v;
	wire v_w5345_v;
	wire v_w6093_v;
	wire v_w6232_v;
	wire v_w1877_v;
	wire v_w4251_v;
	wire v_w6288_v;
	wire v_w4961_v;
	wire v_w7504_v;
	wire v_w7318_v;
	wire v_w1750_v;
	wire v_w5192_v;
	reg v_s254_v;
	wire v_w5279_v;
	wire v_w3294_v;
	wire v_w2990_v;
	wire v_w7910_v;
	wire v_w6782_v;
	wire v_w7914_v;
	wire v_w1797_v;
	wire v_w906_v;
	wire v_w897_v;
	wire v_w172_v;
	wire v_w2739_v;
	wire v_w6947_v;
	wire v_w2330_v;
	wire v_w2861_v;
	wire v_w2987_v;
	wire v_w4299_v;
	wire v_w2768_v;
	wire v_w1026_v;
	wire v_w6856_v;
	wire v_w987_v;
	wire v_w6178_v;
	wire v_w721_v;
	wire v_w7247_v;
	wire v_w2736_v;
	wire v_w7563_v;
	wire v_w7367_v;
	wire v_w1265_v;
	wire v_w249_v;
	wire v_w1600_v;
	wire v_w5292_v;
	wire v_w1584_v;
	wire v_w1980_v;
	wire v_w860_v;
	wire v_w4645_v;
	wire v_w5208_v;
	wire v_w1783_v;
	wire v_w827_v;
	wire v_w8205_v;
	wire v_w3852_v;
	wire v_w7106_v;
	wire v_w5592_v;
	wire v_w7439_v;
	wire v_w1172_v;
	wire v_w3473_v;
	wire v_w339_v;
	wire v_w5918_v;
	wire v_w49_v;
	wire v_w5543_v;
	wire v_w3450_v;
	wire v_w4329_v;
	wire v_w726_v;
	wire v_w7990_v;
	reg v_s179_v;
	wire v_w7001_v;
	wire v_w6391_v;
	wire v_w7010_v;
	wire v_w3589_v;
	wire v_w1891_v;
	wire v_w231_v;
	wire v_w4476_v;
	wire v_w3759_v;
	wire v_w4466_v;
	wire v_w1121_v;
	wire v_w3185_v;
	wire v_w6243_v;
	wire v_w962_v;
	wire v_w3982_v;
	wire v_w5010_v;
	wire v_w1531_v;
	wire v_w1499_v;
	wire v_w4568_v;
	wire v_w4119_v;
	wire v_w3868_v;
	wire v_w6796_v;
	wire v_w922_v;
	wire v_w752_v;
	wire v_w6515_v;
	wire v_w6127_v;
	wire v_w999_v;
	wire v_w6706_v;
	wire v_w1046_v;
	wire v_w4437_v;
	wire v_w5984_v;
	reg v_s151_v;
	wire v_w3785_v;
	wire v_w119_v;
	wire v_w1935_v;
	wire v_w7716_v;
	wire v_w368_v;
	wire v_w6555_v;
	wire v_w1027_v;
	wire v_w7693_v;
	wire v_w6665_v;
	wire v_w6692_v;
	wire v_w87_v;
	wire v_w3947_v;
	wire v_w6602_v;
	wire v_w5819_v;
	wire v_w5542_v;
	wire v_w4619_v;
	wire v_w7278_v;
	wire v_w4806_v;
	wire v_w7008_v;
	wire v_w3507_v;
	wire v_w2197_v;
	wire v_w2170_v;
	wire v_w4362_v;
	wire v_w8099_v;
	wire v_w4174_v;
	wire v_w3411_v;
	wire v_w1723_v;
	wire v_w2994_v;
	wire v_w7895_v;
	wire v_w6176_v;
	wire v_w2613_v;
	wire v_w704_v;
	wire v_w4849_v;
	reg v_s327_v;
	wire v_w498_v;
	wire v_w5680_v;
	wire v_w3100_v;
	wire v_w1650_v;
	wire v_w7796_v;
	wire v_w6126_v;
	wire v_w1805_v;
	wire v_w3973_v;
	wire v_w5337_v;
	wire v_w4044_v;
	wire v_w5886_v;
	wire v_w447_v;
	wire v_w2310_v;
	wire v_w6035_v;
	wire v_w7710_v;
	wire v_w5313_v;
	wire v_w3027_v;
	reg v_s196_v;
	wire v_w5185_v;
	wire v_w875_v;
	wire v_w4688_v;
	wire v_w3718_v;
	reg v_s130_v;
	wire v_w4810_v;
	wire v_w106_v;
	wire v_w146_v;
	wire v_w2527_v;
	wire v_w6139_v;
	wire v_w6607_v;
	wire v_w7401_v;
	wire v_w7629_v;
	wire v_w6273_v;
	wire v_w1358_v;
	wire v_w1166_v;
	reg v_s189_v;
	wire v_w1949_v;
	wire v_w6853_v;
	wire v_w2650_v;
	wire v_w2686_v;
	wire v_w1285_v;
	wire v_w364_v;
	wire v_w2372_v;
	wire v_w1146_v;
	wire v_w5859_v;
	wire v_w3811_v;
	wire v_w1872_v;
	wire v_w6713_v;
	wire v_w1814_v;
	wire v_w7847_v;
	reg v_s407_v;
	wire v_w93_v;
	wire v_w2533_v;
	wire v_w6186_v;
	wire v_w4759_v;
	wire v_w2837_v;
	wire v_w2618_v;
	wire v_w5384_v;
	wire v_w4987_v;
	wire v_w6516_v;
	wire v_w5761_v;
	wire v_w5095_v;
	wire v_w6664_v;
	wire v_w5614_v;
	wire v_w2028_v;
	wire v_w6866_v;
	wire v_w4659_v;
	wire v_w7426_v;
	wire v_w7242_v;
	wire v_w1180_v;
	wire v_w1190_v;
	wire v_w5627_v;
	wire v_w6224_v;
	wire v_w1050_v;
	wire v_w7109_v;
	wire v_w887_v;
	wire v_w1321_v;
	wire v_w4219_v;
	wire v_w2214_v;
	wire v_w6590_v;
	reg v_s346_v;
	wire v_w8026_v;
	reg v_s216_v;
	wire v_w2207_v;
	wire v_w1044_v;
	wire v_w7485_v;
	wire v_w426_v;
	wire v_w6240_v;
	wire v_w377_v;
	wire v_w41_v;
	wire v_w865_v;
	wire v_w5033_v;
	wire v_w6023_v;
	wire v_w589_v;
	wire v_w6765_v;
	wire v_w7930_v;
	wire v_w5156_v;
	wire v_w3339_v;
	wire v_w190_v;
	wire v_w4018_v;
	wire v_w8104_v;
	wire v_w4518_v;
	wire v_w1448_v;
	wire v_w3859_v;
	wire v_w3482_v;
	wire v_w2453_v;
	wire v_w3114_v;
	wire v_w1977_v;
	wire v_w2863_v;
	wire v_w4229_v;
	reg v_s213_v;
	wire v_w4587_v;
	wire v_w1211_v;
	wire v_w7638_v;
	wire v_w337_v;
	wire v_w7600_v;
	wire v_w7231_v;
	wire v_w5722_v;
	wire v_w2673_v;
	wire v_w2190_v;
	wire v_w1571_v;
	wire v_w8043_v;
	wire v_w2081_v;
	wire v_w4710_v;
	wire v_w6345_v;
	wire v_w597_v;
	wire v_w1322_v;
	wire v_w4233_v;
	reg v_s302_v;
	wire v_w2965_v;
	wire v_w4382_v;
	wire v_w8193_v;
	wire v_w357_v;
	wire v_w3862_v;
	wire v_w489_v;
	wire v_w5740_v;
	wire v_w4183_v;
	wire v_w8250_v;
	wire v_w248_v;
	reg v_s397_v;
	wire v_w6081_v;
	wire v_w914_v;
	wire v_w3515_v;
	wire v_w2644_v;
	wire v_w1618_v;
	wire v_w112_v;
	wire v_w6977_v;
	wire v_w3374_v;
	wire v_w6637_v;
	wire v_w7550_v;
	wire v_w5978_v;
	wire v_w1621_v;
	wire v_w4167_v;
	wire v_w5355_v;
	wire v_w2838_v;
	wire v_w6634_v;
	wire v_w5951_v;
	wire v_w4721_v;
	wire v_w3486_v;
	wire v_w581_v;
	wire v_w1947_v;
	wire v_w7507_v;
	wire v_w338_v;
	wire v_w2459_v;
	reg v_s47_v;
	wire v_w1055_v;
	wire v_w1834_v;
	reg v_s518_v;
	wire v_w5231_v;
	wire v_w3068_v;
	wire v_w2221_v;
	wire v_w2286_v;
	wire v_w7976_v;
	reg v_s4_v;
	wire v_w6182_v;
	wire v_w2258_v;
	reg v_s156_v;
	wire v_w3544_v;
	wire v_w5344_v;
	wire v_w3931_v;
	wire v_w4190_v;
	wire v_w3964_v;
	wire v_w2598_v;
	wire v_w4285_v;
	wire v_w4163_v;
	wire v_w5243_v;
	wire v_w3438_v;
	wire v_w4050_v;
	wire v_w2353_v;
	wire v_w2901_v;
	wire v_w6466_v;
	wire v_w1186_v;
	wire v_w6301_v;
	wire v_w5506_v;
	wire v_w3425_v;
	wire v_w4332_v;
	wire v_w8080_v;
	wire v_w1065_v;
	reg v_s292_v;
	wire v_w2440_v;
	wire v_w3750_v;
	wire v_w2021_v;
	reg v_s413_v;
	wire v_w5263_v;
	wire v_w5171_v;
	wire v_w4913_v;
	wire v_w3194_v;
	wire v_w7540_v;
	wire v_w6231_v;
	wire v_w6550_v;
	wire v_w1284_v;
	wire v_w7353_v;
	wire v_w8037_v;
	wire v_w7861_v;
	wire v_w5687_v;
	wire v_w1796_v;
	wire v_w1787_v;
	wire v_w7202_v;
	wire v_w5829_v;
	wire v_w4350_v;
	wire v_w5350_v;
	wire v_w2301_v;
	wire v_w176_v;
	wire v_w2385_v;
	wire v_w7326_v;
	wire v_w5605_v;
	wire v_w767_v;
	wire v_w3963_v;
	wire v_w7314_v;
	wire v_w4266_v;
	wire v_w5781_v;
	wire v_w8009_v;
	wire v_w7265_v;
	wire v_w7103_v;
	reg v_s336_v;
	wire v_w1809_v;
	wire v_w7719_v;
	wire v_w7324_v;
	wire v_w3085_v;
	wire v_w1383_v;
	wire v_w2103_v;
	reg v_s183_v;
	wire v_w7944_v;
	wire v_w5137_v;
	wire v_w1596_v;
	wire v_w7486_v;
	wire v_w771_v;
	wire v_w4714_v;
	wire v_w4327_v;
	wire v_w1323_v;
	wire v_w660_v;
	wire v_w5333_v;
	wire v_w668_v;
	wire v_w821_v;
	wire v_w6776_v;
	wire v_w2836_v;
	wire v_w1899_v;
	wire v_w6161_v;
	wire v_w1173_v;
	wire v_w2007_v;
	wire v_w7235_v;
	wire v_w1656_v;
	wire v_w3072_v;
	wire v_w2433_v;
	wire v_w1687_v;
	wire v_w3330_v;
	wire v_w1806_v;
	wire v_w7203_v;
	wire v_w1998_v;
	wire v_w7089_v;
	wire v_w6669_v;
	wire v_w6254_v;
	wire v_w4128_v;
	wire v_w4585_v;
	wire v_w7270_v;
	wire v_w5166_v;
	wire v_w2556_v;
	reg v_s513_v;
	wire v_w7571_v;
	wire v_w4342_v;
	wire v_w4353_v;
	wire v_w6501_v;
	wire v_w2851_v;
	wire v_w8035_v;
	wire v_w1619_v;
	wire v_w5162_v;
	wire v_w6274_v;
	wire v_w7967_v;
	wire v_w3684_v;
	wire v_w6958_v;
	wire v_w8042_v;
	wire v_w8082_v;
	wire v_w6169_v;
	wire v_w1939_v;
	wire v_w634_v;
	wire v_w5045_v;
	wire v_w4663_v;
	wire v_w3108_v;
	wire v_w5692_v;
	wire v_w2780_v;
	wire v_w4002_v;
	wire v_w2955_v;
	wire v_w7245_v;
	wire v_w6215_v;
	wire v_w1401_v;
	wire v_w7473_v;
	wire v_w8105_v;
	wire v_w1372_v;
	wire v_w7992_v;
	wire v_w3219_v;
	wire v_w5373_v;
	wire v_w1365_v;
	wire v_w537_v;
	wire v_o3_v;
	wire v_w148_v;
	wire v_w7148_v;
	wire v_w5921_v;
	wire v_w6318_v;
	wire v_w2908_v;
	wire v_w1975_v;
	wire v_w4757_v;
	wire v_w354_v;
	wire v_w3535_v;
	wire v_w7299_v;
	wire v_w7892_v;
	wire v_w3783_v;
	wire v_w1849_v;
	wire v_w5123_v;
	wire v_w3427_v;
	wire v_w573_v;
	wire v_w6321_v;
	wire v_w5460_v;
	wire v_w4779_v;
	wire v_w826_v;
	wire v_w1607_v;
	wire v_w4041_v;
	wire v_w873_v;
	wire v_w4686_v;
	wire v_w329_v;
	wire v_w2119_v;
	wire v_w2174_v;
	wire v_w3677_v;
	wire v_w2642_v;
	wire v_w3772_v;
	wire v_w2587_v;
	wire v_w1457_v;
	wire v_w7328_v;
	wire v_w4336_v;
	wire v_w7766_v;
	wire v_w2130_v;
	wire v_w6292_v;
	wire v_w8133_v;
	wire v_w2114_v;
	wire v_w2495_v;
	wire v_w3315_v;
	wire v_w706_v;
	wire v_w1430_v;
	wire v_w5454_v;
	wire v_w3377_v;
	wire v_w3807_v;
	wire v_w5079_v;
	wire v_w7085_v;
	wire v_w5861_v;
	wire v_w5330_v;
	wire v_w1361_v;
	reg v_s451_v;
	wire v_w2608_v;
	wire v_w3882_v;
	wire v_w75_v;
	wire v_w3467_v;
	wire v_w3268_v;
	wire v_w7672_v;
	wire v_w885_v;
	wire v_w5952_v;
	wire v_w107_v;
	wire v_w5521_v;
	wire v_w5088_v;
	wire v_w5556_v;
	wire v_w4897_v;
	wire v_w695_v;
	wire v_w5361_v;
	wire v_w5038_v;
	wire v_w3880_v;
	wire v_w724_v;
	wire v_w1136_v;
	wire v_w909_v;
	wire v_w4904_v;
	reg v_s145_v;
	wire v_w2974_v;
	wire v_w1602_v;
	wire v_w6968_v;
	wire v_w4214_v;
	wire v_w2749_v;
	wire v_w6939_v;
	wire v_w7192_v;
	wire v_o12_v;
	wire v_w5576_v;
	wire v_w6472_v;
	wire v_w7262_v;
	wire v_w3422_v;
	wire v_w1458_v;
	wire v_w2080_v;
	wire v_w3902_v;
	wire v_w1153_v;
	wire v_w6576_v;
	wire v_w3412_v;
	wire v_w7511_v;
	wire v_w7543_v;
	wire v_w749_v;
	wire v_w7298_v;
	wire v_w5034_v;
	wire v_w5367_v;
	wire v_w4578_v;
	wire v_w6386_v;
	wire v_w1832_v;
	wire v_w3514_v;
	wire v_w8238_v;
	wire v_w6026_v;
	wire v_w5520_v;
	wire v_w1090_v;
	wire v_w3092_v;
	wire v_w3707_v;
	wire v_w3351_v;
	wire v_w8050_v;
	wire v_w4094_v;
	wire v_w6614_v;
	wire v_w5256_v;
	wire v_w5046_v;
	wire v_w6068_v;
	wire v_w673_v;
	wire v_w2351_v;
	wire v_w7081_v;
	wire v_w1482_v;
	wire v_w5823_v;
	reg v_s149_v;
	wire v_w6220_v;
	wire v_w4818_v;
	reg v_s334_v;
	wire v_w413_v;
	wire v_w4632_v;
	wire v_w3802_v;
	wire v_w6203_v;
	wire v_w1714_v;
	wire v_w4789_v;
	wire v_w5528_v;
	reg v_s17_v;
	wire v_w682_v;
	wire v_w3537_v;
	wire v_w6506_v;
	wire v_w5306_v;
	wire v_w6786_v;
	reg v_s190_v;
	wire v_w114_v;
	wire v_w98_v;
	wire v_w5679_v;
	wire v_w1756_v;
	wire v_w407_v;
	wire v_w7977_v;
	wire v_w4672_v;
	wire v_w3795_v;
	wire v_w2785_v;
	wire v_w7051_v;
	wire v_w6936_v;
	wire v_w3200_v;
	wire v_w3558_v;
	wire v_w5626_v;
	wire v_w1566_v;
	wire v_w356_v;
	wire v_w655_v;
	wire v_w6821_v;
	wire v_w812_v;
	wire v_w69_v;
	wire v_w5037_v;
	wire v_w2977_v;
	reg v_s398_v;
	wire v_w187_v;
	wire v_w2476_v;
	wire v_w3209_v;
	wire v_w6413_v;
	wire v_w8064_v;
	wire v_w510_v;
	wire v_w861_v;
	wire v_w849_v;
	wire v_w3395_v;
	wire v_w7931_v;
	wire v_w4615_v;
	wire v_w1308_v;
	wire v_w7969_v;
	wire v_w5225_v;
	reg v_s442_v;
	wire v_w3172_v;
	wire v_w1695_v;
	wire v_w6013_v;
	wire v_w6370_v;
	wire v_w3371_v;
	wire v_w609_v;
	wire v_w2743_v;
	wire v_w7558_v;
	wire v_w3661_v;
	wire v_w1962_v;
	wire v_w3937_v;
	wire v_w8032_v;
	wire v_o6_v;
	wire v_w6465_v;
	wire v_w6191_v;
	wire v_w5957_v;
	wire v_w2911_v;
	wire v_w3163_v;
	wire v_w4561_v;
	wire v_w5565_v;
	wire v_w839_v;
	wire v_w2222_v;
	wire v_w5301_v;
	wire v_w3690_v;
	wire v_w4553_v;
	wire v_w3900_v;
	wire v_w85_v;
	wire v_w57_v;
	wire v_w3006_v;
	reg v_s348_v;
	reg v_s419_v;
	wire v_w4257_v;
	wire v_w5135_v;
	wire v_w7189_v;
	wire v_w3403_v;
	wire v_w1219_v;
	reg v_s60_v;
	wire v_w2032_v;
	wire v_w2549_v;
	wire v_w1389_v;
	wire v_w8153_v;
	wire v_w1825_v;
	wire v_w4637_v;
	wire v_w2821_v;
	wire v_w1581_v;
	wire v_w2685_v;
	wire v_w6305_v;
	wire v_w4419_v;
	wire v_w858_v;
	wire v_w2365_v;
	wire v_w4832_v;
	wire v_w3580_v;
	wire v_w2355_v;
	reg v_s232_v;
	reg v_s210_v;
	wire v_w566_v;
	wire v_w854_v;
	wire v_w1079_v;
	wire v_w6034_v;
	wire v_w6327_v;
	wire v_w6142_v;
	wire v_w5828_v;
	wire v_w7791_v;
	wire v_w7276_v;
	wire v_w4760_v;
	reg v_s198_v;
	wire v_w92_v;
	wire v_w3575_v;
	wire v_w7463_v;
	wire v_w1655_v;
	wire v_w2063_v;
	wire v_w7378_v;
	wire v_w3836_v;
	wire v_w6047_v;
	wire v_w7670_v;
	wire v_w1721_v;
	wire v_w5335_v;
	wire v_w2952_v;
	wire v_w2416_v;
	wire v_w4073_v;
	wire v_w3597_v;
	wire v_w269_v;
	wire v_w4724_v;
	wire v_w1390_v;
	wire v_w3634_v;
	wire v_w6025_v;
	wire v_w3773_v;
	wire v_w905_v;
	wire v_w1972_v;
	wire v_w918_v;
	wire v_w3000_v;
	wire v_w8033_v;
	wire v_w6708_v;
	reg v_s120_v;
	wire v_w6247_v;
	reg v_s470_v;
	wire v_w2439_v;
	wire v_w5056_v;
	wire v_o20_v;
	wire v_w2574_v;
	wire v_w7359_v;
	wire v_w7788_v;
	wire v_w6373_v;
	wire v_w1272_v;
	wire v_w572_v;
	wire v_w518_v;
	wire v_w355_v;
	wire v_w3924_v;
	wire v_w3883_v;
	wire v_w222_v;
	wire v_w2256_v;
	wire v_w2012_v;
	wire v_w2361_v;
	wire v_w2260_v;
	wire v_w5120_v;
	wire v_w5158_v;
	reg v_s95_v;
	wire v_w4673_v;
	wire v_w5752_v;
	wire v_w4993_v;
	wire v_w4301_v;
	wire v_w4265_v;
	wire v_w2082_v;
	wire v_w3987_v;
	wire v_w5503_v;
	wire v_w2078_v;
	wire v_w1752_v;
	wire v_w588_v;
	wire v_w3850_v;
	wire v_w3789_v;
	wire v_w2631_v;
	wire v_w7091_v;
	wire v_w212_v;
	wire v_w2726_v;
	wire v_w4872_v;
	wire v_w4652_v;
	wire v_w3766_v;
	wire v_w1717_v;
	wire v_w6352_v;
	wire v_w5360_v;
	wire v_w3423_v;
	wire v_w6748_v;
	wire v_w7315_v;
	wire v_w561_v;
	wire v_w972_v;
	wire v_w1368_v;
	wire v_w4621_v;
	wire v_w3856_v;
	wire v_w3778_v;
	wire v_w6494_v;
	wire v_w4893_v;
	wire v_w1098_v;
	wire v_w2538_v;
	wire v_w1491_v;
	wire v_w1114_v;
	wire v_w6150_v;
	wire v_w1816_v;
	wire v_w5872_v;
	wire v_w2487_v;
	wire v_w331_v;
	wire v_w2057_v;
	wire v_w3060_v;
	wire v_w5494_v;
	wire v_w1413_v;
	wire v_w3673_v;
	wire v_w3010_v;
	reg v_s392_v;
	wire v_w6430_v;
	reg v_s521_v;
	wire v_w3266_v;
	wire v_w2916_v;
	wire v_w4231_v;
	wire v_w3316_v;
	wire v_w4514_v;
	wire v_w312_v;
	wire v_w3096_v;
	wire v_w7214_v;
	wire v_w5741_v;
	wire v_w177_v;
	wire v_w5143_v;
	wire v_w964_v;
	wire v_w5449_v;
	wire v_w1093_v;
	wire v_w3304_v;
	wire v_w7400_v;
	wire v_w2942_v;
	wire v_w3593_v;
	wire v_w72_v;
	wire v_w2591_v;
	wire v_w6668_v;
	wire v_w3075_v;
	wire v_w1248_v;
	wire v_w6140_v;
	wire v_w6088_v;
	wire v_w6635_v;
	wire v_w6629_v;
	wire v_w4985_v;
	wire v_w3504_v;
	wire v_w1928_v;
	wire v_w6175_v;
	wire v_w4863_v;
	wire v_w3817_v;
	wire v_w2253_v;
	wire v_w5787_v;
	reg v_s439_v;
	wire v_w223_v;
	reg v_s264_v;
	wire v_w6451_v;
	wire v_w6064_v;
	wire v_w3969_v;
	wire v_w6617_v;
	wire v_w1638_v;
	wire v_w154_v;
	wire v_w4412_v;
	wire v_w2978_v;
	wire v_w7154_v;
	wire v_w55_v;
	wire v_w257_v;
	wire v_w6193_v;
	reg v_s150_v;
	wire v_w4022_v;
	wire v_w3708_v;
	wire v_w4132_v;
	wire v_w7821_v;
	wire v_w7534_v;
	wire v_w4014_v;
	wire v_w4159_v;
	wire v_w4151_v;
	wire v_w3113_v;
	wire v_w7414_v;
	wire v_w3278_v;
	wire v_w6406_v;
	wire v_w6725_v;
	wire v_w3054_v;
	wire v_w5657_v;
	wire v_w5358_v;
	wire v_w2040_v;
	wire v_w4569_v;
	wire v_w2283_v;
	wire v_w6010_v;
	wire v_w1589_v;
	wire v_w4774_v;
	reg v_s494_v;
	wire v_w5042_v;
	wire v_w2274_v;
	wire v_w4273_v;
	wire v_w990_v;
	wire v_w4200_v;
	wire v_w2751_v;
	wire v_w5862_v;
	wire v_w5069_v;
	wire v_w7646_v;
	wire v_w5003_v;
	wire v_w3333_v;
	wire v_w1301_v;
	wire v_w8132_v;
	wire v_w2501_v;
	wire v_w7206_v;
	wire v_w1506_v;
	wire v_w1889_v;
	wire v_w5409_v;
	wire v_w1486_v;
	wire v_w543_v;
	wire v_w7281_v;
	wire v_w5461_v;
	wire v_w3596_v;
	wire v_w2412_v;
	wire v_w8114_v;
	wire v_w4820_v;
	wire v_w3983_v;
	wire v_w1209_v;
	wire v_w5888_v;
	wire v_w6785_v;
	wire v_w5707_v;
	wire v_w4603_v;
	wire v_w940_v;
	wire v_w7393_v;
	wire v_w6001_v;
	wire v_w4300_v;
	wire v_w6426_v;
	wire v_w5387_v;
	wire v_w8176_v;
	wire v_w2609_v;
	wire v_w1952_v;
	wire v_w3082_v;
	wire v_w5349_v;
	wire v_w8252_v;
	wire v_w5552_v;
	reg v_s349_v;
	wire v_w4976_v;
	wire v_w4630_v;
	wire v_w6310_v;
	wire v_w7440_v;
	wire v_w2299_v;
	wire v_w6536_v;
	wire v_w7963_v;
	wire v_w255_v;
	wire v_w1907_v;
	wire v_w7918_v;
	wire v_w7917_v;
	wire v_w1279_v;
	wire v_w1906_v;
	wire v_w6800_v;
	wire v_w2865_v;
	wire v_w3418_v;
	wire v_w4298_v;
	wire v_w7924_v;
	wire v_w3623_v;
	wire v_w1467_v;
	wire v_w8236_v;
	wire v_w1012_v;
	wire v_w2833_v;
	wire v_w2706_v;
	wire v_w6565_v;
	wire v_w6349_v;
	wire v_w5939_v;
	wire v_w614_v;
	wire v_w7564_v;
	reg v_s236_v;
	wire v_w4815_v;
	wire v_w7417_v;
	wire v_w5774_v;
	wire v_w5673_v;
	wire v_w859_v;
	wire v_w5993_v;
	wire v_w3776_v;
	wire v_w957_v;
	wire v_w7908_v;
	wire v_w8147_v;
	wire v_w646_v;
	wire v_w2641_v;
	wire v_w6572_v;
	wire v_w7019_v;
	wire v_w1314_v;
	wire v_w155_v;
	wire v_w2467_v;
	wire v_w1990_v;
	wire v_w1668_v;
	wire v_w677_v;
	wire v_w5299_v;
	wire v_w2480_v;
	wire v_w4984_v;
	wire v_w6826_v;
	wire v_w6354_v;
	wire v_w2395_v;
	wire v_w6437_v;
	wire v_w1689_v;
	wire v_w2568_v;
	wire v_w1982_v;
	wire v_w3921_v;
	wire v_w5832_v;
	reg v_s54_v;
	wire v_w5533_v;
	wire v_w4660_v;
	wire v_w7734_v;
	wire v_w4302_v;
	wire v_w7213_v;
	wire v_w2061_v;
	wire v_w3483_v;
	wire v_w2651_v;
	wire v_w1103_v;
	wire v_w7301_v;
	wire v_w804_v;
	wire v_w3050_v;
	wire v_w7764_v;
	wire v_w2744_v;
	wire v_w6987_v;
	reg v_s191_v;
	wire v_w5152_v;
	wire v_w7854_v;
	wire v_w478_v;
	wire v_w7530_v;
	wire v_w2101_v;
	wire v_w5709_v;
	wire v_w3408_v;
	wire v_w5611_v;
	wire v_w1699_v;
	wire v_w3716_v;
	wire v_w5570_v;
	wire v_w2907_v;
	wire v_w3282_v;
	wire v_w711_v;
	wire v_w5011_v;
	wire v_w202_v;
	wire v_w2624_v;
	wire v_w7031_v;
	wire v_w5519_v;
	wire v_w1731_v;
	wire v_w104_v;
	wire v_w3162_v;
	wire v_w3289_v;
	wire v_w6770_v;
	wire v_w1979_v;
	wire v_w5773_v;
	wire v_w4503_v;
	wire v_w1405_v;
	wire v_w3324_v;
	wire v_w670_v;
	wire v_w6953_v;
	reg v_s431_v;
	wire v_w3735_v;
	wire v_w7111_v;
	wire v_w5931_v;
	wire v_w768_v;
	reg v_s42_v;
	wire v_w2003_v;
	wire v_w71_v;
	wire v_w5760_v;
	wire v_w3038_v;
	wire v_w37_v;
	wire v_w2731_v;
	wire v_w2213_v;
	wire v_w2975_v;
	wire v_w3616_v;
	wire v_w6498_v;
	wire v_w7210_v;
	wire v_w7628_v;
	wire v_w3576_v;
	wire v_w4577_v;
	wire v_w4722_v;
	wire v_w5738_v;
	wire v_w809_v;
	wire v_w2719_v;
	wire v_w392_v;
	reg v_s353_v;
	wire v_w2868_v;
	wire v_w4508_v;
	wire v_w138_v;
	wire v_w2807_v;
	wire v_w6810_v;
	wire v_w4054_v;
	wire v_w7707_v;
	wire v_w7087_v;
	wire v_w2582_v;
	reg v_s396_v;
	wire v_w2906_v;
	wire v_w2128_v;
	wire v_w2115_v;
	wire v_w6089_v;
	wire v_w2567_v;
	wire v_w3078_v;
	wire v_w2884_v;
	wire v_w7555_v;
	wire v_w5147_v;
	wire v_w2014_v;
	wire v_w1177_v;
	wire v_w2573_v;
	wire v_w5022_v;
	reg v_s437_v;
	wire v_w225_v;
	wire v_w1704_v;
	wire v_w5876_v;
	wire v_w6823_v;
	wire v_w8053_v;
	wire v_w7039_v;
	wire v_w743_v;
	wire v_w7801_v;
	wire v_w1769_v;
	wire v_w3149_v;
	wire v_w3336_v;
	wire v_w644_v;
	wire v_w5919_v;
	wire v_w4478_v;
	wire v_w7120_v;
	wire v_w6615_v;
	wire v_w2323_v;
	wire v_w4982_v;
	wire v_w4402_v;
	wire v_w1645_v;
	wire v_w3323_v;
	reg v_s211_v;
	wire v_w4145_v;
	wire v_w4072_v;
	wire v_w4978_v;
	wire v_w5343_v;
	wire v_w8054_v;
	wire v_w1534_v;
	wire v_w3586_v;
	wire v_w7070_v;
	wire v_w5435_v;
	wire v_w8199_v;
	wire v_w1340_v;
	wire v_w6286_v;
	reg v_s71_v;
	wire v_w3801_v;
	wire v_w3540_v;
	wire v_w7184_v;
	wire v_w5535_v;
	wire v_w722_v;
	wire v_w4080_v;
	wire v_w5402_v;
	wire v_w4047_v;
	wire v_w2292_v;
	wire v_w3872_v;
	wire v_w7599_v;
	wire v_w2311_v;
	wire v_w2919_v;
	wire v_w786_v;
	wire v_w4967_v;
	wire v_w937_v;
	wire v_w6510_v;
	wire v_w1074_v;
	wire v_w2514_v;
	wire v_w3794_v;
	wire v_w3925_v;
	wire v_w5845_v;
	reg v_s408_v;
	wire v_w6523_v;
	wire v_w4004_v;
	wire v_w3117_v;
	wire v_w1514_v;
	wire v_w168_v;
	wire v_w2238_v;
	wire v_w2475_v;
	wire v_w7394_v;
	wire v_w3146_v;
	wire v_w7040_v;
	wire v_w4243_v;
	wire v_w1002_v;
	wire v_w302_v;
	wire v_w4137_v;
	wire v_w1056_v;
	wire v_w1052_v;
	wire v_w4060_v;
	wire v_w3198_v;
	wire v_w5468_v;
	wire v_w7146_v;
	wire v_w4258_v;
	wire v_w6038_v;
	wire v_w5516_v;
	reg v_s269_v;
	wire v_w4479_v;
	wire v_w5155_v;
	wire v_w3737_v;
	wire v_w7509_v;
	wire v_w6385_v;
	wire v_w982_v;
	wire v_w3934_v;
	wire v_w6598_v;
	wire v_w7985_v;
	wire v_w927_v;
	wire v_w4328_v;
	wire v_w6238_v;
	wire v_w3112_v;
	reg v_s194_v;
	wire v_w4246_v;
	wire v_w1878_v;
	reg v_s275_v;
	wire v_w5000_v;
	wire v_w1230_v;
	wire v_w2463_v;
	wire v_w3837_v;
	wire v_w7946_v;
	wire v_w6690_v;
	wire v_w8117_v;
	wire v_w7937_v;
	wire v_w4153_v;
	wire v_w6022_v;
	wire v_w3134_v;
	wire v_w2947_v;
	wire v_w2243_v;
	wire v_w4009_v;
	wire v_w3258_v;
	wire v_w5163_v;
	wire v_w5332_v;
	wire v_w6961_v;
	wire v_w3009_v;
	wire v_w6869_v;
	wire v_w3474_v;
	wire v_w4361_v;
	wire v_w5265_v;
	wire v_w4783_v;
	wire v_w4711_v;
	wire v_w7130_v;
	wire v_w3142_v;
	wire v_w4185_v;
	wire v_w4098_v;
	wire v_w4717_v;
	wire v_w4017_v;
	wire v_w8187_v;
	wire v_w6375_v;
	reg v_s182_v;
	wire v_w6894_v;
	wire v_w5757_v;
	wire v_w3188_v;
	wire v_w5639_v;
	wire v_w4846_v;
	wire v_w3044_v;
	wire v_w1631_v;
	wire v_w6179_v;
	wire v_w2347_v;
	wire v_w4590_v;
	wire v_w1586_v;
	wire v_w4108_v;
	wire v_w985_v;
	wire v_w1738_v;
	wire v_w4683_v;
	wire v_w1813_v;
	wire v_w2909_v;
	wire v_w4385_v;
	wire v_w943_v;
	wire v_w4234_v;
	wire v_w4370_v;
	wire v_w4821_v;
	wire v_w8213_v;
	reg v_s245_v;
	wire v_w1268_v;
	wire v_w5447_v;
	wire v_w6219_v;
	wire v_o9_v;
	wire v_w3320_v;
	wire v_w4012_v;
	wire v_w1895_v;
	wire v_w5696_v;
	wire v_w7531_v;
	wire v_w3274_v;
	wire v_w5814_v;
	reg v_s499_v;
	wire v_w89_v;
	wire v_w7551_v;
	wire v_w97_v;
	wire v_w7500_v;
	wire v_w4924_v;
	wire v_w1651_v;
	wire v_w3915_v;
	wire v_w7252_v;
	wire v_w5180_v;
	wire v_w6079_v;
	wire v_w4541_v;
	wire v_o21_v;
	wire v_w4411_v;
	wire v_w1520_v;
	wire v_w7277_v;
	wire v_w2005_v;
	reg v_s365_v;
	wire v_w3091_v;
	wire v_w7399_v;
	wire v_w7312_v;
	wire v_w3813_v;
	wire v_w6100_v;
	wire v_w301_v;
	wire v_w7887_v;
	wire v_w3547_v;
	wire v_w7323_v;
	wire v_w4983_v;
	wire v_w6030_v;
	wire v_w7916_v;
	wire v_w6724_v;
	wire v_w1815_v;
	wire v_w198_v;
	wire v_w514_v;
	wire v_w3758_v;
	wire v_w2205_v;
	wire v_w5363_v;
	wire v_w7413_v;
	wire v_w5950_v;
	wire v_w1360_v;
	wire v_w5836_v;
	wire v_w7375_v;
	reg v_s489_v;
	wire v_w129_v;
	wire v_w6969_v;
	wire v_w6144_v;
	wire v_w406_v;
	wire v_w6133_v;
	wire v_w659_v;
	wire v_w267_v;
	wire v_w515_v;
	wire v_w7090_v;
	wire v_w5525_v;
	wire v_w2619_v;
	wire v_w6228_v;
	wire v_w5812_v;
	wire v_w7102_v;
	wire v_w6798_v;
	wire v_w577_v;
	wire v_w825_v;
	wire v_w4142_v;
	wire v_w6149_v;
	wire v_w5177_v;
	wire v_w6265_v;
	wire v_w116_v;
	wire v_w3065_v;
	wire v_w3835_v;
	wire v_w2870_v;
	wire v_w5669_v;
	wire v_w6087_v;
	wire v_w3087_v;
	wire v_w3954_v;
	wire v_w6951_v;
	wire v_w6008_v;
	wire v_w6648_v;
	wire v_w1910_v;
	wire v_w5550_v;
	wire v_w5161_v;
	wire v_w1352_v;
	reg v_s280_v;
	wire v_w1551_v;
	wire v_w1240_v;
	wire v_w4359_v;
	wire v_w6449_v;
	wire v_w4441_v;
	reg v_s256_v;
	wire v_w7445_v;
	wire v_w1880_v;
	wire v_w5703_v;
	wire v_w5379_v;
	wire v_w5668_v;
	wire v_w5972_v;
	wire v_w3555_v;
	wire v_w5414_v;
	wire v_w8188_v;
	wire v_w791_v;
	wire v_w3356_v;
	wire v_w871_v;
	wire v_w2657_v;
	wire v_w965_v;
	wire v_w2235_v;
	reg v_s447_v;
	reg v_s261_v;
	wire v_w5025_v;
	wire v_w2455_v;
	wire v_w2096_v;
	reg v_s127_v;
	wire v_w1319_v;
	wire v_w528_v;
	wire v_w2006_v;
	wire v_w5587_v;
	wire v_w1614_v;
	reg v_s2_v;
	wire v_w7297_v;
	wire v_w7855_v;
	wire v_w8012_v;
	wire v_w5544_v;
	reg v_s27_v;
	wire v_w380_v;
	wire v_w855_v;
	wire v_w617_v;
	wire v_w7038_v;
	wire v_w3641_v;
	wire v_w3181_v;
	wire v_w345_v;
	wire v_w6261_v;
	wire v_w6431_v;
	wire v_w1548_v;
	wire v_w621_v;
	wire v_w3792_v;
	wire v_w3256_v;
	wire v_w7319_v;
	wire v_w7283_v;
	wire v_w2180_v;
	wire v_w6441_v;
	wire v_w5151_v;
	wire v_w6138_v;
	reg v_s11_v;
	reg v_s147_v;
	reg v_s281_v;
	wire v_w6212_v;
	wire v_w6984_v;
	wire v_w5061_v;
	wire v_w8116_v;
	wire v_w2989_v;
	wire v_w974_v;
	wire v_w599_v;
	wire v_w237_v;
	wire v_w7411_v;
	wire v_w7215_v;
	wire v_w5254_v;
	wire v_w7117_v;
	wire v_w516_v;
	wire v_w4850_v;
	wire v_w6207_v;
	wire v_w340_v;
	wire v_w636_v;
	wire v_w3686_v;
	wire v_w416_v;
	wire v_w2715_v;
	wire v_w3671_v;
	wire v_w2411_v;
	wire v_w2281_v;
	wire v_w744_v;
	wire v_w3445_v;
	wire v_w2603_v;
	wire v_w4464_v;
	wire v_w5218_v;
	wire v_w6971_v;
	wire v_w1088_v;
	wire v_w3036_v;
	wire v_w3024_v;
	wire v_w2371_v;
	wire v_w3165_v;
	wire v_w6408_v;
	wire v_w4684_v;
	reg v_s93_v;
	wire v_w5716_v;
	wire v_w1031_v;
	wire v_w5489_v;
	wire v_w5127_v;
	wire v_w2985_v;
	wire v_w280_v;
	wire v_w2322_v;
	wire v_w3290_v;
	wire v_w6925_v;
	wire v_w1123_v;
	wire v_w3700_v;
	wire v_w479_v;
	wire v_w2778_v;
	wire v_w1329_v;
	wire v_o10_v;
	wire v_w7999_v;
	wire v_w7780_v;
	wire v_w1781_v;
	wire v_w2380_v;
	reg v_s383_v;
	wire v_w3157_v;
	wire v_w669_v;
	wire v_w1119_v;
	wire v_w6799_v;
	wire v_w3846_v;
	wire v_w1840_v;
	wire v_w3610_v;
	wire v_w6673_v;
	wire v_w6448_v;
	wire v_w234_v;
	wire v_w676_v;
	wire v_w233_v;
	wire v_w4146_v;
	wire v_w799_v;
	wire v_w633_v;
	wire v_w2633_v;
	reg v_s126_v;
	wire v_w4888_v;
	wire v_w5370_v;
	wire v_w7795_v;
	wire v_w1451_v;
	wire v_w4870_v;
	reg v_s153_v;
	wire v_w7163_v;
	reg v_s128_v;
	wire v_w158_v;
	wire v_w197_v;
	wire v_w5539_v;
	wire v_w5159_v;
	wire v_w6793_v;
	wire v_w6923_v;
	wire v_w7641_v;
	reg v_s330_v;
	wire v_w8189_v;
	wire v_w5851_v;
	wire v_w2734_v;
	wire v_w1269_v;
	wire v_w951_v;
	wire v_w3424_v;
	wire v_w6416_v;
	wire v_w1916_v;
	wire v_w7129_v;
	wire v_w6121_v;
	wire v_w6571_v;
	reg v_s293_v;
	wire v_w3663_v;
	wire v_w7781_v;
	wire v_w4805_v;
	wire v_w6541_v;
	wire v_w6102_v;
	wire v_w5144_v;
	reg v_s108_v;
	wire v_w6880_v;
	reg v_s177_v;
	wire v_w3747_v;
	wire v_w3041_v;
	wire v_w5662_v;
	wire v_w4900_v;
	wire v_w1644_v;
	wire v_w7617_v;
	wire v_w2891_v;
	reg v_s277_v;
	wire v_w3675_v;
	wire v_w7835_v;
	wire v_w4495_v;
	wire v_w1927_v;
	wire v_w7360_v;
	wire v_w2389_v;
	reg v_s289_v;
	wire v_w4197_v;
	wire v_w7140_v;
	wire v_w998_v;
	reg v_s415_v;
	wire v_w2179_v;
	wire v_w1684_v;
	wire v_w3806_v;
	wire v_w2635_v;
	wire v_w5153_v;
	wire v_w7173_v;
	wire v_w1135_v;
	wire v_w7024_v;
	wire v_w3654_v;
	wire v_w4109_v;
	wire v_w7698_v;
	wire v_w4554_v;
	wire v_w4371_v;
	wire v_w6905_v;
	wire v_w3440_v;
	wire v_w5269_v;
	wire v_w67_v;
	reg v_s515_v;
	wire v_w4039_v;
	wire v_w2569_v;
	wire v_w6753_v;
	wire v_w6582_v;
	wire v_w2840_v;
	wire v_w4333_v;
	wire v_w3436_v;
	wire v_w7819_v;
	wire v_w5002_v;
	wire v_w6214_v;
	wire v_w7982_v;
	wire v_w2451_v;
	wire v_w3125_v;
	wire v_w2133_v;
	wire v_w1696_v;
	wire v_w8154_v;
	wire v_w6780_v;
	wire v_w5028_v;
	wire v_w2674_v;
	wire v_w4745_v;
	wire v_w4946_v;
	wire v_w5769_v;
	wire v_w6152_v;
	wire v_w1951_v;
	wire v_w2553_v;
	wire v_w3106_v;
	wire v_w4100_v;
	wire v_w4038_v;
	wire v_w3975_v;
	reg v_s509_v;
	wire v_w6409_v;
	wire v_w7836_v;
	wire v_w5086_v;
	wire v_w6945_v;
	wire v_w2161_v;
	wire v_w5712_v;
	wire v_w446_v;
	reg v_s22_v;
	wire v_w1345_v;
	wire v_w5820_v;
	reg v_s514_v;
	wire v_o11_v;
	wire v_w7107_v;
	wire v_w6289_v;
	wire v_w7723_v;
	wire v_w4097_v;
	reg v_s462_v;
	wire v_w3167_v;
	reg v_s250_v;
	wire v_w4928_v;
	wire v_w2147_v;
	wire v_w6353_v;
	wire v_w2991_v;
	wire v_w384_v;
	wire v_w4963_v;
	wire v_w1822_v;
	wire v_w4248_v;
	wire v_w6603_v;
	wire v_w1305_v;
	wire v_w2009_v;
	wire v_w4051_v;
	wire v_w3475_v;
	reg v_s343_v;
	wire v_w7650_v;
	wire v_w7524_v;
	wire v_w8149_v;
	wire v_w6258_v;
	wire v_w5327_v;
	wire v_w6057_v;
	wire v_w1118_v;
	reg v_s10_v;
	wire v_w31_v;
	wire v_w8088_v;
	wire v_w61_v;
	wire v_w6339_v;
	wire v_w2442_v;
	wire v_w5786_v;
	wire v_w6410_v;
	wire v_w2124_v;
	wire v_w1399_v;
	wire v_w7320_v;
	wire v_w6694_v;
	wire v_w6535_v;
	wire v_w2472_v;
	wire v_w4618_v;
	wire v_w5366_v;
	wire v_w3302_v;
	wire v_w5685_v;
	wire v_w4700_v;
	wire v_w3285_v;
	wire v_w4641_v;
	wire v_w5223_v;
	wire v_w6661_v;
	wire v_w418_v;
	wire v_w7496_v;
	wire v_w1158_v;
	wire v_w1789_v;
	wire v_w5107_v;
	wire v_w200_v;
	wire v_w2002_v;
	wire v_w5179_v;
	wire v_w7651_v;
	wire v_w313_v;
	wire v_w6729_v;
	wire v_w6389_v;
	wire v_w244_v;
	wire v_w2710_v;
	wire v_w2928_v;
	wire v_w2341_v;
	wire v_w6056_v;
	wire v_w2626_v;
	wire v_w5695_v;
	wire v_w896_v;
	wire v_w1083_v;
	wire v_w51_v;
	reg v_s352_v;
	wire v_w7002_v;
	wire v_w7282_v;
	wire v_w7625_v;
	wire v_w1475_v;
	wire v_w2008_v;
	wire v_w6046_v;
	wire v_w3692_v;
	wire v_w3_v;
	wire v_w3236_v;
	wire v_w6778_v;
	wire v_w2498_v;
	wire v_w5247_v;
	wire v_w485_v;
	wire v_w4565_v;
	wire v_w6718_v;
	wire v_w2273_v;
	wire v_w1477_v;
	wire v_w7833_v;
	wire v_w102_v;
	wire v_w4894_v;
	wire v_w303_v;
	wire v_w7480_v;
	wire v_w6118_v;
	wire v_w7219_v;
	wire v_w3015_v;
	wire v_w3141_v;
	wire v_w911_v;
	wire v_w1449_v;
	reg v_s123_v;
	wire v_w5008_v;
	wire v_w8221_v;
	wire v_w7110_v;
	wire v_w5122_v;
	wire v_w4838_v;
	wire v_w1522_v;
	wire v_w7922_v;
	wire v_w389_v;
	wire v_w4980_v;
	wire v_w246_v;
	wire v_w807_v;
	wire v_w8228_v;
	wire v_w2803_v;
	wire v_w6364_v;
	wire v_w6312_v;
	reg v_s443_v;
	wire v_w4260_v;
	wire v_w3935_v;
	wire v_w427_v;
	wire v_w4392_v;
	wire v_w6048_v;
	wire v_w6671_v;
	wire v_w5675_v;
	wire v_w6732_v;
	wire v_w1495_v;
	wire v_w6787_v;
	wire v_w862_v;
	wire v_w981_v;
	wire v_w6279_v;
	wire v_w2210_v;
	reg v_s344_v;
	wire v_w3032_v;
	wire v_w6839_v;
	wire v_w7454_v;
	wire v_w5255_v;
	wire v_w2386_v;
	wire v_w7499_v;
	wire v_w2388_v;
	wire v_w7479_v;
	wire v_w6870_v;
	wire v_o8_v;
	wire v_w7702_v;
	wire v_w4292_v;
	wire v_w546_v;
	wire v_w5172_v;
	wire v_w3484_v;
	wire v_w3414_v;
	wire v_w5746_v;
	reg v_s418_v;
	wire v_w6707_v;
	wire v_w5524_v;
	wire v_w210_v;
	wire v_w3284_v;
	wire v_w5678_v;
	wire v_w3410_v;
	wire v_w6728_v;
	wire v_w1973_v;
	wire v_w3843_v;
	wire v_w1503_v;
	wire v_w2391_v;
	wire v_w6137_v;
	wire v_w5380_v;
	wire v_w1630_v;
	wire v_w2167_v;
	wire v_w1524_v;
	wire v_w2031_v;
	wire v_w7424_v;
	wire v_w1022_v;
	wire v_w6343_v;
	wire v_w147_v;
	wire v_w5138_v;
	wire v_w7288_v;
	wire v_w746_v;
	wire v_w5148_v;
	wire v_w1157_v;
	wire v_w2141_v;
	wire v_w118_v;
	wire v_w2934_v;
	wire v_w3489_v;
	wire v_w7475_v;
	wire v_w1893_v;
	wire v_w1582_v;
	wire v_w3855_v;
	wire v_w4695_v;
	wire v_w7978_v;
	wire v_w5501_v;
	wire v_w5253_v;
	wire v_w5420_v;
	wire v_w5251_v;
	wire v_w3966_v;
	wire v_w7305_v;
	wire v_w5227_v;
	wire v_w6225_v;
	wire v_w6382_v;
	wire v_w7438_v;
	wire v_w28_v;
	wire v_w5963_v;
	wire v_w893_v;
	wire v_w330_v;
	wire v_w3088_v;
	wire v_w5681_v;
	wire v_w2931_v;
	wire v_w973_v;
	wire v_w3025_v;
	reg v_s215_v;
	wire v_w5300_v;
	wire v_w7906_v;
	wire v_w2236_v;
	wire v_w7776_v;
	wire v_w4454_v;
	wire v_w1422_v;
	wire v_w462_v;
	wire v_w7349_v;
	wire v_w7952_v;
	wire v_w4713_v;
	wire v_w7921_v;
	wire v_w7878_v;
	wire v_w4462_v;
	wire v_w3711_v;
	wire v_w5964_v;
	wire v_w5369_v;
	wire v_w6851_v;
	wire v_w2027_v;
	wire v_w5507_v;
	wire v_w1215_v;
	wire v_w3511_v;
	wire v_w5425_v;
	wire v_w2554_v;
	wire v_w5099_v;
	wire v_w1014_v;
	wire v_w3048_v;
	wire v_w124_v;
	wire v_w1976_v;
	reg v_s90_v;
	wire v_w8101_v;
	wire v_w3699_v;
	wire v_w3821_v;
	wire v_w2168_v;
	wire v_w2497_v;
	wire v_w2324_v;
	wire v_w7510_v;
	wire v_w5372_v;
	wire v_w7212_v;
	wire v_w4186_v;
	wire v_w3881_v;
	wire v_w7965_v;
	wire v_w7652_v;
	wire v_w1971_v;
	wire v_w6067_v;
	wire v_w953_v;
	wire v_w2026_v;
	wire v_w7841_v;
	wire v_w7879_v;
	wire v_w4129_v;
	wire v_w4348_v;
	wire v_w5968_v;
	wire v_w5866_v;
	reg v_s433_v;
	wire v_w6942_v;
	wire v_w2334_v;
	wire v_w605_v;
	wire v_w7669_v;
	wire v_w7062_v;
	wire v_w8230_v;
	wire v_w4738_v;
	wire v_w1444_v;
	wire v_w22_v;
	wire v_w2656_v;
	wire v_w2072_v;
	wire v_w3203_v;
	wire v_w8074_v;
	wire v_w6970_v;
	wire v_w3592_v;
	wire v_w494_v;
	wire v_w4032_v;
	wire v_w6890_v;
	wire v_w6532_v;
	wire v_w5749_v;
	wire v_w1423_v;
	wire v_w3938_v;
	wire v_o7_v;
	wire v_w1017_v;
	wire v_w1334_v;
	wire v_w789_v;
	wire v_w335_v;
	wire v_w7108_v;
	wire v_w3746_v;
	wire v_w3170_v;
	wire v_w1111_v;
	wire v_w3174_v;
	wire v_w798_v;
	wire v_w5314_v;
	wire v_w5636_v;
	wire v_w4892_v;
	wire v_w8046_v;
	wire v_w4782_v;
	wire v_w4278_v;
	wire v_w1035_v;
	reg v_s410_v;
	wire v_w5326_v;
	wire v_w4939_v;
	wire v_w3159_v;
	wire v_w5960_v;
	wire v_w471_v;
	wire v_w863_v;
	wire v_w3460_v;
	wire v_w5858_v;
	wire v_w1327_v;
	wire v_w2469_v;
	wire v_w165_v;
	wire v_w295_v;
	wire v_w8068_v;
	wire v_w1433_v;
	wire v_w4028_v;
	wire v_w955_v;
	wire v_w8124_v;
	wire v_w8130_v;
	wire v_w5618_v;
	wire v_w7630_v;
	wire v_w2319_v;
	wire v_w4859_v;
	wire v_w2444_v;
	wire v_w1421_v;
	wire v_w8025_v;
	wire v_w7139_v;
	wire v_w2376_v;
	wire v_w3842_v;
	wire v_w1080_v;
	wire v_w4655_v;
	wire v_w6929_v;
	wire v_w6016_v;
	wire v_w833_v;
	wire v_w1216_v;
	wire v_w6401_v;
	wire v_w63_v;
	wire v_w4702_v;
	wire v_w5413_v;
	wire v_w2596_v;
	wire v_w1623_v;
	wire v_w1957_v;
	wire v_w6857_v;
	wire v_w1521_v;
	wire v_w7150_v;
	wire v_w3917_v;
	wire v_w5512_v;
	wire v_w774_v;
	wire v_w3840_v;
	wire v_w2348_v;
	wire v_w742_v;
	wire v_w8168_v;
	reg v_s323_v;
	wire v_w1249_v;
	wire v_w3179_v;
	wire v_w5174_v;
	wire v_w1604_v;
	wire v_w4058_v;
	wire v_w4422_v;
	wire v_w7434_v;
	wire v_w2971_v;
	wire v_w6508_v;
	wire v_w2912_v;
	wire v_w5383_v;
	wire v_w503_v;
	wire v_w5509_v;
	wire v_w134_v;
	wire v_w7464_v;
	wire v_w5329_v;
	reg v_s221_v;
	wire v_w8107_v;
	wire v_w3516_v;
	wire v_w5076_v;
	wire v_w1373_v;
	wire v_w5339_v;
	wire v_w2502_v;
	wire v_w691_v;
	wire v_w5775_v;
	wire v_w2079_v;
	wire v_w3808_v;
	wire v_w7046_v;
	wire v_w7042_v;
	wire v_w6313_v;
	wire v_w5453_v;
	wire v_w3107_v;
	wire v_w2873_v;
	wire v_w6306_v;
	wire v_w3896_v;
	wire v_w6222_v;
	wire v_w6517_v;
	wire v_w1425_v;
	reg v_s485_v;
	wire v_w1094_v;
	wire v_w6817_v;
	wire v_w167_v;
	wire v_w7455_v;
	wire v_w6907_v;
	wire v_w4640_v;
	wire v_w1547_v;
	wire v_w1311_v;
	wire v_w1363_v;
	wire v_w6721_v;
	wire v_w3977_v;
	wire v_w2446_v;
	wire v_w4903_v;
	wire v_w1068_v;
	wire v_w6824_v;
	wire v_w1539_v;
	wire v_w5486_v;
	wire v_w8067_v;
	wire v_w2799_v;
	wire v_w7626_v;
	wire v_w7420_v;
	wire v_w252_v;
	wire v_w592_v;
	wire v_w360_v;
	wire v_w7736_v;
	wire v_w3669_v;
	wire v_w501_v;
	reg v_s482_v;
	wire v_w7158_v;
	wire v_w46_v;
	wire v_w5282_v;
	reg v_s235_v;
	wire v_w6471_v;
	reg v_s26_v;
	wire v_w4534_v;
	wire v_w5765_v;
	wire v_w4509_v;
	wire v_w7831_v;
	wire v_w2151_v;
	wire v_w6085_v;
	wire v_w8140_v;
	wire v_w2278_v;
	wire v_w7444_v;
	wire v_w4491_v;
	wire v_w3725_v;
	wire v_w1393_v;
	wire v_w6077_v;
	wire v_w1597_v;
	wire v_w5903_v;
	wire v_w1406_v;
	wire v_w4520_v;
	wire v_w1845_v;
	wire v_w584_v;
	wire v_w4428_v;
	wire v_w1622_v;
	wire v_w3150_v;
	wire v_w7696_v;
	wire v_w5597_v;
	wire v_w1149_v;
	wire v_w5428_v;
	wire v_w3992_v;
	wire v_w2721_v;
	wire v_w1370_v;
	wire v_w497_v;
	wire v_w1817_v;
	wire v_w3697_v;
	wire v_w6886_v;
	wire v_w7025_v;
	wire v_w4612_v;
	wire v_w7181_v;
	wire v_w8109_v;
	wire v_w4232_v;
	wire v_w6050_v;
	wire v_w7246_v;
	wire v_w2466_v;
	wire v_w4791_v;
	wire v_w1603_v;
	wire v_w567_v;
	wire v_w5538_v;
	wire v_w3497_v;
	wire v_w490_v;
	wire v_w2589_v;
	wire v_w6336_v;
	wire v_w3246_v;
	wire v_w7284_v;
	wire v_w1875_v;
	wire v_w2212_v;
	wire v_w5839_v;
	wire v_w2252_v;
	wire v_w7186_v;
	wire v_w320_v;
	wire v_w7957_v;
	wire v_w2401_v;
	wire v_w2699_v;
	wire v_w2571_v;
	wire v_w2824_v;
	wire v_w6827_v;
	wire v_w1400_v;
	wire v_w2270_v;
	wire v_w3124_v;
	wire v_w6876_v;
	wire v_w6993_v;
	wire v_w540_v;
	wire v_w2593_v;
	wire v_w6360_v;
	wire v_w640_v;
	wire v_w6542_v;
	wire v_w3600_v;
	wire v_w3439_v;
	wire v_w2452_v;
	wire v_w6014_v;
	wire v_w4741_v;
	wire v_w7639_v;
	wire v_w3228_v;
	wire v_w7566_v;
	wire v_w4160_v;
	reg v_s299_v;
	wire v_w2832_v;
	wire v_w3858_v;
	wire v_w1986_v;
	wire v_w5566_v;
	wire v_w7757_v;
	wire v_w7296_v;
	wire v_w8020_v;
	wire v_w5569_v;
	wire v_w433_v;
	wire v_w7354_v;
	wire v_w3352_v;
	wire v_w3223_v;
	wire v_w3121_v;
	wire v_w1316_v;
	wire v_w6256_v;
	wire v_w2183_v;
	wire v_w2927_v;
	wire v_w627_v;
	wire v_w444_v;
	wire v_w4268_v;
	wire v_w1011_v;
	wire v_w5994_v;
	wire v_w1690_v;
	wire v_w5296_v;
	wire v_w595_v;
	wire v_w95_v;
	wire v_w1049_v;
	wire v_w2271_v;
	wire v_w7345_v;
	wire v_w7559_v;
	wire v_w4293_v;
	wire v_w73_v;
	reg v_s152_v;
	wire v_w2615_v;
	wire v_w4836_v;
	wire v_w4776_v;
	wire v_w2015_v;
	wire v_w1530_v;
	wire v_w2765_v;
	wire v_w8004_v;
	wire v_w5388_v;
	wire v_w5633_v;
	wire v_w7826_v;
	reg v_s88_v;
	wire v_w6719_v;
	wire v_w6356_v;
	reg v_s55_v;
	reg v_s137_v;
	wire v_w3153_v;
	wire v_w7223_v;
	wire v_w6234_v;
	wire v_w2586_v;
	reg v_s432_v;
	wire v_w7361_v;
	wire v_w2646_v;
	wire v_w4207_v;
	wire v_w1904_v;
	wire v_w2383_v;
	wire v_w748_v;
	wire v_w50_v;
	wire v_w2137_v;
	wire v_w1808_v;
	wire v_w4873_v;
	wire v_w3510_v;
	wire v_w3672_v;
	wire v_w5572_v;
	wire v_w3341_v;
	wire v_w5068_v;
	wire v_w1874_v;
	wire v_w8249_v;
	reg v_s163_v;
	wire v_w1671_v;
	wire v_w3061_v;
	wire v_w1161_v;
	wire v_w1516_v;
	wire v_w5087_v;
	reg v_s92_v;
	wire v_w7830_v;
	wire v_w8162_v;
	wire v_w6599_v;
	wire v_w7790_v;
	reg v_s136_v;
	wire v_w6838_v;
	wire v_w7190_v;
	wire v_w5979_v;
	wire v_w171_v;
	wire v_w810_v;
	wire v_w6727_v;
	wire v_w4935_v;
	wire v_w2224_v;
	wire v_w8158_v;
	wire v_w7269_v;
	wire v_w4010_v;
	reg v_s291_v;
	wire v_w6066_v;
	wire v_w3035_v;
	wire v_w6006_v;
	wire v_w2899_v;
	wire v_w2264_v;
	wire v_w8040_v;
	wire v_w7981_v;
	wire v_w683_v;
	wire v_w2481_v;
	wire v_w6759_v;
	wire v_w1469_v;
	wire v_w2234_v;
	wire v_w2964_v;
	wire v_w4034_v;
	wire v_w4937_v;
	wire v_w3139_v;
	wire v_w256_v;
	wire v_w3461_v;
	wire v_w1929_v;
	wire v_w126_v;
	wire v_w5091_v;
	reg v_s464_v;
	wire v_w3825_v;
	reg v_s197_v;
	wire v_w3744_v;
	wire v_w414_v;
	wire v_w6505_v;
	wire v_w4066_v;
	wire v_w3144_v;
	wire v_w3827_v;
	wire v_w7653_v;
	wire v_w2941_v;
	reg v_s510_v;
	wire v_w3218_v;
	wire v_w6333_v;
	wire v_w6054_v;
	wire v_w7017_v;
	wire v_o5_v;
	wire v_w79_v;
	wire v_w2810_v;
	wire v_w1855_v;
	wire v_w7994_v;
	wire v_w7497_v;
	wire v_w6687_v;
	wire v_w2512_v;
	wire v_w2173_v;
	wire v_w2622_v;
	wire v_w2374_v;
	wire v_w2869_v;
	wire v_w6656_v;
	wire v_w1568_v;
	wire v_w4720_v;
	wire v_w4908_v;
	wire v_w6746_v;
	wire v_w2443_v;
	reg v_s516_v;
	wire v_w692_v;
	reg v_s227_v;
	wire v_w4857_v;
	wire v_w4715_v;
	wire v_w729_v;
	wire v_w2419_v;
	wire v_w4896_v;
	wire v_w3039_v;
	wire v_w6659_v;
	wire v_w1351_v;
	wire v_w2428_v;
	wire v_w3476_v;
	wire v_w6973_v;
	wire v_w5232_v;
	wire v_w2249_v;
	wire v_w476_v;
	wire v_w8049_v;
	wire v_w6553_v;
	reg v_s340_v;
	wire v_w4092_v;
	wire v_w6552_v;
	wire v_w2515_v;
	wire v_w3328_v;
	wire v_w2152_v;
	wire v_w5316_v;
	wire v_w7508_v;
	wire v_w1758_v;
	wire v_w1476_v;
	wire v_w4796_v;
	wire v_w5244_v;
	wire v_w1921_v;
	wire v_w3740_v;
	wire v_w7421_v;
	wire v_w4964_v;
	wire v_w7166_v;
	wire v_w3479_v;
	wire v_w6924_v;
	wire v_w3748_v;
	reg v_s288_v;
	wire v_w6745_v;
	wire v_w4571_v;
	wire v_w2425_v;
	wire v_w6893_v;
	wire v_w4456_v;
	wire v_w3135_v;
	wire v_w4029_v;
	wire v_w4530_v;
	wire v_w371_v;
	reg v_s169_v;
	wire v_w1698_v;
	wire v_w5191_v;
	wire v_w4706_v;
	wire v_w1434_v;
	wire v_w7182_v;
	wire v_w3689_v;
	wire v_w565_v;
	wire v_w533_v;
	wire v_w5949_v;
	wire v_w4440_v;
	wire v_w4662_v;
	wire v_w6735_v;
	wire v_w2797_v;
	wire v_w1887_v;
	wire v_w2186_v;
	wire v_w5510_v;
	wire v_w1735_v;
	wire v_w7679_v;
	wire v_w448_v;
	wire v_w3175_v;
	wire v_w6842_v;
	wire v_w7582_v;
	wire v_w2774_v;
	wire v_w3448_v;
	wire v_w4202_v;
	wire v_w3536_v;
	wire v_w4778_v;
	wire v_w7815_v;
	wire v_w2143_v;
	wire v_w5856_v;
	wire v_w7634_v;
	reg v_s9_v;
	wire v_w7837_v;
	wire v_w1288_v;
	reg v_s129_v;
	wire v_w959_v;
	wire v_w1102_v;
	wire v_w7726_v;
	wire v_w8203_v;
	reg v_s51_v;
	wire v_w6445_v;
	wire v_w5459_v;
	wire v_w4910_v;
	wire v_w5288_v;
	wire v_w1407_v;
	wire v_w5097_v;
	wire v_w4264_v;
	wire v_w6462_v;
	reg v_s412_v;
	reg v_s324_v;
	wire v_w7643_v;
	wire v_w5271_v;
	wire v_w8234_v;
	wire v_w3379_v;
	wire v_w513_v;
	wire v_w3939_v;
	wire v_w5312_v;
	wire v_w7239_v;
	reg v_s477_v;
	wire v_w8094_v;
	wire v_w2513_v;
	wire v_w4215_v;
	wire v_w2695_v;
	wire v_w1143_v;
	wire v_w2545_v;
	wire v_w3469_v;
	wire v_w1198_v;
	wire v_w2740_v;
	wire v_w3962_v;
	wire v_w1356_v;
	wire v_w2782_v;
	wire v_w2060_v;
	wire v_w4600_v;
	wire v_w7968_v;
	wire v_w3090_v;
	wire v_w5809_v;
	reg v_s283_v;
	wire v_w6895_v;
	wire v_w5956_v;
	wire v_w6803_v;
	wire v_w7183_v;
	wire v_w4226_v;
	wire v_w5936_v;
	wire v_w3989_v;
	wire v_w3612_v;
	wire v_w8163_v;
	wire v_w7852_v;
	wire v_w2075_v;
	reg v_s382_v;
	wire v_w3155_v;
	wire v_w8021_v;
	wire v_w290_v;
	wire v_w6537_v;
	wire v_w3583_v;
	wire v_w1384_v;
	wire v_w14_v;
	wire v_w2688_v;
	reg v_s411_v;
	wire v_w2069_v;
	wire v_w7149_v;
	wire v_w7381_v;
	wire v_w1201_v;
	wire v_w6108_v;
	wire v_w6367_v;
	wire v_w7126_v;
	wire v_w4055_v;
	wire v_w7704_v;
	wire v_w346_v;
	wire v_w3283_v;
	wire v_w3211_v;
	wire v_w7885_v;
	wire v_w6877_v;
	wire v_w3204_v;
	wire v_w755_v;
	wire v_w5248_v;
	wire v_w7539_v;
	wire v_w2730_v;
	wire v_w449_v;
	wire v_w3086_v;
	wire v_w3653_v;
	wire v_w5081_v;
	wire v_w2516_v;
	wire v_w1772_v;
	wire v_w5200_v;
	wire v_w6253_v;
	wire v_w4560_v;
	wire v_w3847_v;
	wire v_w1106_v;
	wire v_w7218_v;
	wire v_w5113_v;
	wire v_w5057_v;
	wire v_w7261_v;
	wire v_w2572_v;
	wire v_w3694_v;
	wire v_w6158_v;
	wire v_w1130_v;
	wire v_w2566_v;
	wire v_w3224_v;
	wire v_w6522_v;
	wire v_w7114_v;
	wire v_w151_v;
	wire v_w7226_v;
	wire v_w5473_v;
	wire v_w5776_v;
	wire v_w396_v;
	wire v_w253_v;
	wire v_w2915_v;
	wire v_w1231_v;
	wire v_w6257_v;
	wire v_w1324_v;
	wire v_w6277_v;
	wire v_w7874_v;
	wire v_w530_v;
	wire v_w4358_v;
	wire v_w1639_v;
	wire v_w1847_v;
	wire v_w2056_v;
	wire v_w7468_v;
	wire v_w6005_v;
	wire v_w1839_v;
	wire v_w1412_v;
	wire v_w6731_v;
	wire v_w3624_v;
	wire v_w2074_v;
	wire v_w4949_v;
	wire v_w4528_v;
	wire v_w2261_v;
	wire v_w1481_v;
	wire v_w1988_v;
	wire v_w7133_v;
	wire v_w6033_v;
	wire v_w4582_v;
	wire v_w5640_v;
	wire v_w7730_v;
	wire v_w7100_v;
	wire v_w6106_v;
	wire v_w1261_v;
	wire v_w7251_v;
	wire v_w594_v;
	wire v_w1724_v;
	wire v_w2561_v;
	wire v_w6366_v;
	wire v_w4453_v;
	wire v_w4962_v;
	wire v_w2628_v;
	wire v_w843_v;
	wire v_w1646_v;
	wire v_w3980_v;
	wire v_w2665_v;
	wire v_w6395_v;
	wire v_w5906_v;
	wire v_w3229_v;
	wire v_w8081_v;
	wire v_w3208_v;
	wire v_w4307_v;
	wire v_w3326_v;
	wire v_w6843_v;
	wire v_w7583_v;
	wire v_w2177_v;
	reg v_s157_v;
	reg v_s325_v;
	wire v_w6705_v;
	wire v_w4562_v;
	wire v_w1033_v;
	wire v_w4956_v;
	wire v_w6828_v;
	wire v_w2897_v;
	wire v_w1515_v;
	wire v_w3667_v;
	wire v_w7607_v;
	wire v_w484_v;
	wire v_w4868_v;
	wire v_w7596_v;
	wire v_w3122_v;
	wire v_w2610_v;
	wire v_w5607_v;
	wire v_w8017_v;
	wire v_w324_v;
	wire v_w4992_v;
	wire v_w1594_v;
	wire v_w7909_v;
	wire v_w400_v;
	wire v_w5444_v;
	wire v_w7157_v;
	wire v_w376_v;
	wire v_w1913_v;
	wire v_w8121_v;
	wire v_w5573_v;
	wire v_w526_v;
	wire v_w6859_v;
	wire v_w4395_v;
	wire v_w1468_v;
	wire v_w7113_v;
	wire v_w1037_v;
	wire v_w7733_v;
	wire v_w7761_v;
	wire v_w8122_v;
	wire v_w4614_v;
	wire v_w2879_v;
	wire v_w3731_v;
	wire v_w2431_v;
	wire v_w394_v;
	wire v_w3115_v;
	wire v_w5285_v;
	wire v_w4693_v;
	wire v_w772_v;
	wire v_w3426_v;
	wire v_w1730_v;
	wire v_w81_v;
	wire v_w4500_v;
	wire v_w5470_v;
	wire v_w8177_v;
	wire v_w828_v;
	wire v_w6200_v;
	reg v_s255_v;
	wire v_w4733_v;
	reg v_s36_v;
	wire v_w4486_v;
	wire v_w1510_v;
	wire v_w2969_v;
	wire v_w1375_v;
	wire v_w7768_v;
	wire v_w2750_v;
	wire v_w6369_v;
	wire v_w2796_v;
	wire v_w2808_v;
	wire v_w4111_v;
	wire v_w3681_v;
	wire v_w3259_v;
	wire v_w7799_v;
	wire v_w2160_v;
	wire v_w7498_v;
	wire v_w5995_v;
	wire v_w199_v;
	wire v_w8172_v;
	wire v_w1004_v;
	wire v_w3265_v;
	wire v_w1295_v;
	wire v_w6909_v;
	wire v_w8223_v;
	wire v_w7119_v;
	wire v_w4981_v;
	wire v_w803_v;
	wire v_w3539_v;
	wire v_w164_v;
	wire v_w6989_v;
	wire v_w6573_v;
	wire v_w6663_v;
	wire v_w6468_v;
	wire v_w4506_v;
	wire v_w3629_v;
	wire v_w68_v;
	reg v_s354_v;
	wire v_w6551_v;
	wire v_w2461_v;
	wire v_w2486_v;
	wire v_w3132_v;
	wire v_w7436_v;
	wire v_w732_v;
	wire v_w1487_v;
	wire v_w1007_v;
	wire v_w1064_v;
	wire v_w5235_v;
	wire v_w3166_v;
	wire v_w6985_v;
	wire v_w1974_v;
	wire v_w8202_v;
	wire v_w1700_v;
	wire v_w511_v;
	wire v_w4844_v;
	wire v_w853_v;
	wire v_w8233_v;
	wire v_w2397_v;
	wire v_w6995_v;
	wire v_w1658_v;
	wire v_w7065_v;
	wire v_w6814_v;
	wire v_w5146_v;
	wire v_w7591_v;
	wire v_w1206_v;
	wire v_w966_v;
	wire v_w3958_v;
	wire v_w3177_v;
	wire v_w3943_v;
	wire v_w7465_v;
	wire v_w1392_v;
	wire v_w6347_v;
	wire v_w4773_v;
	wire v_w6117_v;
	wire v_w582_v;
	wire v_w7026_v;
	wire v_w3638_v;
	wire v_w7487_v;
	wire v_w980_v;
	wire v_w7593_v;
	wire v_w5522_v;
	wire v_w4256_v;
	wire v_w6815_v;
	wire v_w4680_v;
	wire v_w1722_v;
	wire v_w6818_v;
	wire v_w311_v;
	wire v_w4091_v;
	wire v_w4308_v;
	wire v_w4418_v;
	wire v_w8003_v;
	wire v_w90_v;
	wire v_w8215_v;
	wire v_w2599_v;
	wire v_w204_v;
	wire v_w2792_v;
	wire v_w2544_v;
	wire v_w1179_v;
	wire v_w930_v;
	wire v_w115_v;
	wire v_w1152_v;
	reg v_s406_v;
	wire v_w1480_v;
	wire v_w7156_v;
	wire v_w5229_v;
	wire v_w6300_v;
	wire v_w6340_v;
	wire v_w6561_v;
	wire v_w5490_v;
	wire v_w3976_v;
	wire v_w2135_v;
	wire v_w5693_v;
	wire v_w5670_v;
	wire v_w477_v;
	wire v_w731_v;
	wire v_w2288_v;
	wire v_w7597_v;
	wire v_w7427_v;
	wire v_w1233_v;
	wire v_w2847_v;
	wire v_w7482_v;
	reg v_s113_v;
	wire v_w4220_v;
	wire v_w6504_v;
	wire v_w1898_v;
	wire v_w7667_v;
	wire v_w3520_v;
	wire v_w1532_v;
	wire v_w6833_v;
	wire v_w7515_v;
	wire v_w7923_v;
	wire v_w6199_v;
	wire v_w4548_v;
	wire v_w649_v;
	wire v_w7703_v;
	wire v_w1882_v;
	wire v_w123_v;
	wire v_w4690_v;
	wire v_w2083_v;
	wire v_w1385_v;
	wire v_w4668_v;
	wire v_w3069_v;
	wire v_w2317_v;
	wire v_w6992_v;
	wire v_w3604_v;
	wire v_w1330_v;
	wire v_w3552_v;
	wire v_w697_v;
	wire v_w5595_v;
	wire v_w2804_v;
	wire v_w1277_v;
	wire v_w6646_v;
	wire v_w7391_v;
	wire v_w2943_v;
	wire v_w5270_v;
	wire v_w2268_v;
	wire v_w3350_v;
	wire v_w2489_v;
	wire v_w7059_v;
	wire v_w5706_v;
	wire v_w2902_v;
	wire v_w7385_v;
	wire v_w2920_v;
	wire v_w2043_v;
	wire v_w287_v;
	wire v_w1359_v;
	wire v_w6460_v;
	wire v_w6195_v;
	wire v_w740_v;
	wire v_w664_v;
	wire v_w6060_v;
	wire v_w7516_v;
	wire v_w5671_v;
	wire v_w938_v;
	wire v_w5175_v;
	wire v_w4533_v;
	wire v_w910_v;
	wire v_w4812_v;
	wire v_w2275_v;
	wire v_w6962_v;
	wire v_w7101_v;
	wire v_w4646_v;
	wire v_w6875_v;
	wire v_w867_v;
	wire v_w7866_v;
	wire v_w6439_v;
	wire v_w1036_v;
	wire v_w3660_v;
	wire v_w3554_v;
	wire v_w8152_v;
	reg v_s87_v;
	wire v_w1378_v;
	wire v_w7238_v;
	reg v_s474_v;
	wire v_w4296_v;
	wire v_w2693_v;
	wire v_w7838_v;
	wire v_w100_v;
	wire v_w7654_v;
	wire v_w3105_v;
	reg v_s175_v;
	wire v_w4626_v;
	wire v_w4297_v;
	wire v_w7356_v;
	wire v_w1795_v;
	wire v_w1831_v;
	wire v_w4784_v;
	wire v_w8106_v;
	wire v_w7151_v;
	wire v_w3936_v;
	wire v_w5131_v;
	wire v_w5801_v;
	wire v_w7263_v;
	wire v_w3275_v;
	wire v_w2649_v;
	wire v_w7682_v;
	wire v_w4753_v;
	wire v_w7627_v;
	wire v_w5893_v;
	wire v_w4954_v;
	wire v_w2711_v;
	wire v_w284_v;
	wire v_w3066_v;
	wire v_w919_v;
	wire v_w2839_v;
	wire v_w4003_v;
	wire v_w8019_v;
	wire v_w5666_v;
	wire v_w279_v;
	wire v_w8058_v;
	wire v_w1665_v;
	wire v_w7327_v;
	wire v_w7343_v;
	reg v_s205_v;
	wire v_w6278_v;
	wire v_w4950_v;
	wire v_w5534_v;
	wire v_w4769_v;
	wire v_w5643_v;
	reg v_s223_v;
	wire v_w4376_v;
	wire v_w716_v;
	wire v_w1362_v;
	wire v_w4737_v;
	wire v_w2580_v;
	wire v_w3201_v;
	wire v_w5432_v;
	wire v_w2864_v;
	wire v_w1649_v;
	wire v_w3253_v;
	wire v_w6916_v;
	wire v_w3506_v;
	reg v_s103_v;
	wire v_w1633_v;
	wire v_w4239_v;
	wire v_w3509_v;
	wire v_w2632_v;
	wire v_w7688_v;
	wire v_w2944_v;
	reg v_s496_v;
	wire v_w2136_v;
	wire v_w6259_v;
	wire v_w7347_v;
	wire v_w553_v;
	wire v_w6720_v;
	wire v_w1583_v;
	wire v_w1133_v;
	reg v_s371_v;
	wire v_w2312_v;
	wire v_w1948_v;
	wire v_w5424_v;
	wire v_w5199_v;
	wire v_w7061_v;
	wire v_w610_v;
	wire v_w1541_v;
	wire v_w7743_v;
	wire v_w94_v;
	wire v_w2164_v;
	wire v_w4249_v;
	wire v_w5119_v;
	wire v_w2423_v;
	wire v_w6443_v;
	wire v_w1504_v;
	reg v_s390_v;
	wire v_w191_v;
	wire v_w7807_v;
	wire v_w5395_v;
	wire v_w3206_v;
	wire v_w7988_v;
	wire v_w924_v;
	wire v_w5418_v;
	wire v_w4310_v;
	wire v_w568_v;
	wire v_w7785_v;
	wire v_w5331_v;
	wire v_w4414_v;
	wire v_w579_v;
	wire v_w4212_v;
	wire v_w3545_v;
	wire v_w848_v;
	wire v_w6652_v;
	wire v_w229_v;
	wire v_w4915_v;
	wire v_w262_v;
	wire v_w5196_v;
	wire v_w8139_v;
	wire v_w3303_v;
	wire v_w1835_v;
	wire v_w997_v;
	wire v_w4117_v;
	wire v_w1196_v;
	reg v_s206_v;
	wire v_w6685_v;
	wire v_w3472_v;
	wire v_w436_v;
	wire v_w7082_v;
	wire v_w5186_v;
	wire v_o2_v;
	wire v_w8181_v;
	wire v_w2993_v;
	wire v_w892_v;
	wire v_w6358_v;
	wire v_w4502_v;
	wire v_w2215_v;
	wire v_w353_v;
	wire v_w3498_v;
	reg v_s166_v;
	wire v_w2605_v;
	wire v_w3053_v;
	wire v_w20_v;
	reg v_s114_v;
	wire v_w2871_v;
	wire v_w623_v;
	wire v_w7877_v;
	wire v_w690_v;
	wire v_w370_v;
	reg v_s195_v;
	wire v_w2970_v;
	wire v_w3387_v;
	wire v_w7862_v;
	wire v_w1380_v;
	wire v_w4252_v;
	wire v_w2748_v;
	wire v_w8171_v;
	wire v_w1922_v;
	wire v_w4294_v;
	wire v_w5925_v;
	wire v_w1737_v;
	wire v_w6558_v;
	wire v_w7092_v;
	wire v_w6061_v;
	wire v_w2362_v;
	reg v_s290_v;
	wire v_w2790_v;
	wire v_w7886_v;
	wire v_w5321_v;
	wire v_w6633_v;
	wire v_w2961_v;
	wire v_w7377_v;
	wire v_w5149_v;
	wire v_w7657_v;
	wire v_w4801_v;
	wire v_w5054_v;
	wire v_w2979_v;
	wire v_w5021_v;
	wire v_w1267_v;
	wire v_w6474_v;
	wire v_w5750_v;
	wire v_w1298_v;
	wire v_w1335_v;
	wire v_w6107_v;
	wire v_w7175_v;
	reg v_s359_v;
	wire v_w2406_v;
	wire v_w3849_v;
	wire v_w1558_v;
	wire v_w3959_v;
	wire v_w1128_v;
	wire v_w5391_v;
	wire v_w1484_v;
	wire v_w1167_v;
	wire v_w4015_v;
	reg v_s364_v;
	wire v_w2898_v;
	wire v_w7720_v;
	wire v_w3319_v;
	wire v_w6280_v;
	reg v_s49_v;
	wire v_w3417_v;
	wire v_w7991_v;
	reg v_s139_v;
	wire v_w7677_v;
	wire v_w8143_v;
	wire v_w4827_v;
	wire v_w1163_v;
	wire v_w1968_v;
	wire v_w4696_v;
	wire v_w5182_v;
	wire v_w3343_v;
	wire v_w736_v;
	wire v_w2652_v;
	wire v_w2534_v;
	wire v_w5895_v;
	reg v_s282_v;
	wire v_w7514_v;
	wire v_w2393_v;
	wire v_w8113_v;
	wire v_w2779_v;
	wire v_w1901_v;
	wire v_w6852_v;
	wire v_w1280_v;
	wire v_w5206_v;
	wire v_w3532_v;
	reg v_s99_v;
	reg v_s53_v;
	wire v_w4941_v;
	wire v_w3685_v;
	reg v_s414_v;
	wire v_w7987_v;
	wire v_w2818_v;
	reg v_s378_v;
	wire v_w7741_v;
	wire v_w638_v;
	wire v_w2968_v;
	wire v_w5474_v;
	wire v_w1342_v;
	wire v_w6245_v;
	wire v_w3570_v;
	wire v_w6844_v;
	wire v_w2185_v;
	wire v_w6129_v;
	wire v_w7406_v;
	wire v_w5134_v;
	wire v_w4211_v;
	wire v_w7637_v;
	wire v_w7222_v;
	wire v_w1025_v;
	wire v_w6999_v;
	reg v_s203_v;
	wire v_w5280_v;
	wire v_w7752_v;
	reg v_s242_v;
	wire v_w3299_v;
	wire v_w717_v;
	wire v_w8211_v;
	wire v_w3775_v;
	wire v_w2262_v;
	wire v_w7585_v;
	wire v_w4986_v;
	wire v_w4749_v;
	reg v_s154_v;
	wire v_w2611_v;
	wire v_w1303_v;
	wire v_w4572_v;
	wire v_w2559_v;
	wire v_w1127_v;
	wire v_w3331_v;
	wire v_w3787_v;
	wire v_w1403_v;
	wire v_w7389_v;
	wire v_w77_v;
	wire v_w1518_v;
	wire v_w7840_v;
	wire v_w5850_v;
	wire v_w7975_v;
	wire v_w5982_v;
	wire v_w2125_v;
	reg v_s295_v;
	wire v_w3688_v;
	wire v_w4829_v;
	wire v_w2684_v;
	wire v_w5452_v;
	wire v_w5463_v;
	wire v_w5455_v;
	wire v_w3154_v;
	wire v_w1718_v;
	wire v_w4799_v;
	wire v_w5754_v;
	wire v_w4557_v;
	wire v_w1148_v;
	wire v_w1613_v;
	wire v_w3786_v;
	wire v_w1470_v;
	wire v_w8186_v;
	wire v_w6073_v;
	wire v_w4309_v;
	reg v_s91_v;
	wire v_w5588_v;
	wire v_w6374_v;
	reg v_s142_v;
	wire v_w6972_v;
	wire v_w6112_v;
	wire v_w3790_v;
	wire v_w2995_v;
	wire v_w6920_v;
	reg v_s98_v;
	wire v_w3913_v;
	wire v_w7228_v;
	reg v_s466_v;
	wire v_w2938_v;
	wire v_w6837_v;
	wire v_w7760_v;
	wire v_w4316_v;
	wire v_w2036_v;
	wire v_w76_v;
	wire v_w6433_v;
	wire v_w4692_v;
	wire v_w7532_v;
	wire v_w3021_v;
	wire v_w6711_v;
	wire v_w7084_v;
	wire v_w4204_v;
	wire v_w6529_v;
	reg v_s318_v;
	wire v_w4394_v;
	wire v_w8217_v;
	wire v_w8248_v;
	wire v_w4494_v;
	wire v_w6070_v;
	reg v_s212_v;
	wire v_w3774_v;
	wire v_w2729_v;
	wire v_w7236_v;
	wire v_w3368_v;
	wire v_w6601_v;
	wire v_w3784_v;
	wire v_w7256_v;
	wire v_w2066_v;
	wire v_w4882_v;
	wire v_w7339_v;
	wire v_w7993_v;
	wire v_w5986_v;
	wire v_w5909_v;
	wire v_w6262_v;
	wire v_w895_v;
	wire v_w564_v;
	wire v_w2802_v;
	wire v_w247_v;
	wire v_w4628_v;
	reg v_s164_v;
	wire v_w4357_v;
	wire v_w4811_v;
	wire v_w3543_v;
	wire v_w2297_v;
	wire v_w5892_v;
	wire v_w5184_v;
	wire v_w1564_v;
	wire v_w4481_v;
	wire v_w4194_v;
	wire v_w7875_v;
	wire v_w5052_v;
	wire v_w3617_v;
	wire v_w328_v;
	wire v_w6290_v;
	wire v_w2110_v;
	reg v_s486_v;
	wire v_w7519_v;
	wire v_w2298_v;
	wire v_w2788_v;
	wire v_w7372_v;
	wire v_w268_v;
	wire v_w2998_v;
	wire v_w2664_v;
	wire v_w266_v;
	wire v_w1235_v;
	reg v_s326_v;
	wire v_w466_v;
	wire v_w1932_v;
	wire v_w3437_v;
	reg v_s81_v;
	wire v_w6847_v;
	wire v_w5297_v;
	wire v_w2890_v;
	wire v_w3861_v;
	wire v_w8010_v;
	wire v_w3703_v;
	wire v_w4463_v;
	wire v_w5267_v;
	wire v_w6227_v;
	wire v_w7035_v;
	wire v_w432_v;
	wire v_w7407_v;
	wire v_w6604_v;
	wire v_w2350_v;
	wire v_w4447_v;
	wire v_w1076_v;
	wire v_w3234_v;
	wire v_w3782_v;
	wire v_w6415_v;
	wire v_w1632_v;
	wire v_w2427_v;
	wire v_w6883_v;
	wire v_w4306_v;
	wire v_w5181_v;
	wire v_w2812_v;
	wire v_w7774_v;
	wire v_w6263_v;
	wire v_w3390_v;
	wire v_w3369_v;
	wire v_w6610_v;
	wire v_w5755_v;
	wire v_w3161_v;
	wire v_w7545_v;
	wire v_w5574_v;
	wire v_w3345_v;
	wire v_w4599_v;
	wire v_w1920_v;
	reg v_s337_v;
	wire v_w321_v;
	wire v_w558_v;
	wire v_w5249_v;
	wire v_w3585_v;
	wire v_w5701_v;
	wire v_w5511_v;
	wire v_w2450_v;
	wire v_w6213_v;
	wire v_w7174_v;
	wire v_w2178_v;
	wire v_w2318_v;
	wire v_w7045_v;
	wire v_w3191_v;
	wire v_w8013_v;
	wire v_w6493_v;
	wire v_w6211_v;
	wire v_w7581_v;
	reg v_s193_v;
	wire v_w5145_v;
	wire v_w7681_v;
	wire v_w7797_v;
	wire v_w4068_v;
	wire v_w453_v;
	wire v_w1478_v;
	wire v_w1141_v;
	wire v_w4168_v;
	wire v_w7191_v;
	wire v_w8127_v;
	wire v_w6091_v;
	wire v_w3749_v;
	wire v_w5049_v;
	wire v_w2948_v;
	wire v_w96_v;
	wire v_o1_v;
	wire v_w5867_v;
	wire v_w2682_v;
	wire v_w2922_v;
	wire v_w1746_v;
	wire v_w5806_v;
	wire v_w5169_v;
	wire v_w74_v;
	wire v_w1523_v;
	reg v_s370_v;
	wire v_w2625_v;
	wire v_w1994_v;
	wire v_w5485_v;
	wire v_w7005_v;
	reg v_s467_v;
	wire v_w992_v;
	wire v_w5245_v;
	wire v_w580_v;
	reg v_s305_v;
	wire v_w5917_v;
	wire v_w1070_v;
	wire v_w2496_v;
	wire v_w2775_v;
	wire v_w1771_v;
	wire v_w3116_v;
	wire v_w3956_v;
	wire v_w7740_v;
	wire v_w1162_v;
	wire v_w2225_v;
	wire v_w3443_v;
	wire v_w6187_v;
	wire v_w47_v;
	wire v_w7602_v;
	wire v_w2477_v;
	wire v_w7633_v;
	wire v_w412_v;
	wire v_w6533_v;
	wire v_w3370_v;
	reg v_s481_v;
	wire v_w719_v;
	wire v_w6170_v;
	wire v_w7023_v;
	wire v_w297_v;
	reg v_s161_v;
	wire v_w7404_v;
	wire v_w6802_v;
	wire v_w8090_v;
	wire v_w8112_v;
	wire v_w5527_v;
	wire v_w1567_v;
	wire v_w2720_v;
	wire v_w4914_v;
	wire v_w2247_v;
	wire v_w1492_v;
	wire v_w2017_v;
	wire v_w7370_v;
	wire v_w845_v;
	wire v_w6124_v;
	wire v_w7230_v;
	wire v_w1867_v;
	wire v_w1938_v;
	wire v_w3325_v;
	wire v_w1930_v;
	wire v_w2022_v;
	reg v_s140_v;
	wire v_w4093_v;
	wire v_w3026_v;
	wire v_w1533_v;
	wire v_w1833_v;
	wire v_w4965_v;
	wire v_w5217_v;
	wire v_w4973_v;
	wire v_w802_v;
	wire v_w2203_v;
	wire v_w3145_v;
	wire v_w1678_v;
	wire v_w1785_v;
	wire v_w2980_v;
	wire v_w3059_v;
	wire v_w8207_v;
	wire v_w4658_v;
	wire v_w1081_v;
	wire v_w3664_v;
	wire v_w7459_v;
	reg v_s214_v;
	wire v_w1894_v;
	wire v_w5955_v;
	wire v_w7280_v;
	wire v_w8146_v;
	wire v_w2623_v;
	wire v_w7250_v;
	wire v_w8242_v;
	wire v_w2874_v;
	reg v_s278_v;
	wire v_w4597_v;
	wire v_w3019_v;
	wire v_w7396_v;
	wire v_w2309_v;
	wire v_w7680_v;
	wire v_w2420_v;
	wire v_w7379_v;
	wire v_w2030_v;
	reg v_s167_v;
	wire v_w101_v;
	wire v_w889_v;
	reg v_s475_v;
	wire v_w6693_v;
	wire v_w4526_v;
	wire v_w5030_v;
	wire v_w7529_v;
	reg v_s25_v;
	wire v_w7358_v;
	wire v_w6959_v;
	wire v_w4793_v;
	wire v_w5352_v;
	wire v_w1770_v;
	wire v_w1742_v;
	reg v_s28_v;
	wire v_w3195_v;
	wire v_w1200_v;
	wire v_w3531_v;
	wire v_w5495_v;
	wire v_w7227_v;
	wire v_w2875_v;
	wire v_w916_v;
	wire v_w6309_v;
	wire v_w1220_v;
	wire v_w1826_v;
	wire v_w1028_v;
	reg v_s380_v;
	wire v_w4288_v;
	wire v_w3851_v;
	reg v_s367_v;
	wire v_w1885_v;
	wire v_w1544_v;
	wire v_w1803_v;
	wire v_w5777_v;
	wire v_w4344_v;
	wire v_w17_v;
	wire v_w461_v;
	wire v_w5730_v;
	wire v_w7441_v;
	wire v_w3864_v;
	wire v_o22_v;
	wire v_w4694_v;
	wire v_w2787_v;
	wire v_w6205_v;
	wire v_w6754_v;
	wire v_w4379_v;
	wire v_w4529_v;
	wire v_w7588_v;
	wire v_w2370_v;
	wire v_w1748_v;
	wire v_w3503_v;
	wire v_w7642_v;
	wire v_w5213_v;
	reg v_s117_v;
	wire v_w2004_v;
	wire v_w797_v;
	wire v_w1091_v;
	wire v_w7747_v;
	wire v_w215_v;
	wire v_w365_v;
	wire v_w4756_v;
	wire v_w5736_v;
	wire v_w4112_v;
	wire v_w4349_v;
	wire v_w6739_v;
	wire v_w2607_v;
	wire v_w3542_v;
	wire v_w783_v;
	wire v_w6738_v;
	wire v_w7063_v;
	wire v_w3815_v;
	wire v_w7171_v;
	wire v_w7533_v;
	wire v_w7355_v;
	wire v_w3186_v;
	wire v_w1561_v;
	wire v_w557_v;
	wire v_w1527_v;
	wire v_w7180_v;
	wire v_w7934_v;
	wire v_w6597_v;
	wire v_w8241_v;
	wire v_w4922_v;
	wire v_w4101_v;
	wire v_w6435_v;
	wire v_w864_v;
	wire v_w7048_v;
	wire v_w6109_v;
	wire v_w2058_v;
	reg v_s285_v;
	wire v_w3393_v;
	wire v_w6361_v;
	wire v_w5997_v;
	wire v_w7196_v;
	wire v_w6450_v;
	wire v_w2701_v;
	wire v_w3867_v;
	wire v_w7336_v;
	wire v_w4687_v;
	wire v_w2402_v;
	wire v_w5791_v;
	wire v_w3138_v;
	wire v_w6612_v;
	wire v_w7729_v;
	wire v_w221_v;
	wire v_w5371_v;
	wire v_w7904_v;
	wire v_w492_v;
	wire v_w2835_v;
	wire v_w2226_v;
	wire v_w6986_v;
	wire v_w4865_v;
	wire v_w5660_v;
	wire v_w787_v;
	wire v_w5205_v;
	wire v_w7664_v;
	wire v_w7383_v;
	reg v_s355_v;
	wire v_w6194_v;
	wire v_w2460_v;
	wire v_w6294_v;
	wire v_w7408_v;
	wire v_w631_v;
	wire v_w1672_v;
	wire v_w1818_v;
	wire v_w3495_v;
	wire v_w7860_v;
	wire v_o19_v;
	reg v_s116_v;
	wire v_w3084_v;
	wire v_w2896_v;
	wire v_w3603_v;
	reg v_s454_v;
	wire v_w7955_v;
	wire v_w6201_v;
	wire v_w2344_v;
	wire v_w2054_v;
	wire v_w4416_v;
	wire v_w5642_v;
	wire v_w781_v;
	wire v_w2045_v;
	wire v_w5882_v;
	reg v_s294_v;
	wire v_w1234_v;
	wire v_w3622_v;
	wire v_w547_v;
	wire v_w4948_v;
	reg v_s85_v;
	wire v_w1673_v;
	wire v_w7894_v;
	wire v_w6269_v;
	wire v_w1765_v;
	wire v_w2062_v;
	wire v_w2421_v;
	wire v_w8175_v;
	wire v_w3429_v;
	wire v_w6938_v;
	wire v_w4023_v;
	wire v_w7724_v;
	wire v_w836_v;
	wire v_w3841_v;
	wire v_w5864_v;
	wire v_w4189_v;
	wire v_w4401_v;
	wire v_w5407_v;
	wire v_w4007_v;
	reg v_s18_v;
	wire v_w2800_v;
	wire v_w6660_v;
	wire v_w132_v;
	reg v_s30_v;
	wire v_w3739_v;
	wire v_w195_v;
	wire v_w585_v;
	wire v_w5904_v;
	wire v_w230_v;
	wire v_w5029_v;
	wire v_w263_v;
	wire v_w5480_v;
	reg v_s276_v;
	wire v_w5233_v;
	wire v_w4134_v;
	wire v_w3300_v;
	wire v_w3430_v;
	wire v_w6702_v;
	wire v_w2999_v;
	wire v_w1900_v;
	wire v_w2842_v;
	wire v_w288_v;
	wire v_w3594_v;
	wire v_w4669_v;
	reg v_s504_v;
	wire v_w7580_v;
	wire v_w8092_v;
	wire v_w281_v;
	wire v_w3271_v;
	wire v_w5031_v;
	wire v_w745_v;
	wire v_w7488_v;
	wire v_w4409_v;
	wire v_w3521_v;
	wire v_w5891_v;
	wire v_w3464_v;
	wire v_w460_v;
	wire v_w5117_v;
	wire v_w5059_v;
	wire v_w7384_v;
	wire v_w6736_v;
	wire v_w1058_v;
	wire v_w2099_v;
	wire v_w7466_v;
	wire v_w4120_v;
	reg v_s270_v;
	wire v_w3541_v;
	wire v_w1841_v;
	wire v_w5434_v;
	reg v_s100_v;
	wire v_w5913_v;
	wire v_w3242_v;
	wire v_w3866_v;
	wire v_w1820_v;
	wire v_w3465_v;
	wire v_w1409_v;
	wire v_w8220_v;
	wire v_w5_v;
	wire v_w470_v;
	wire v_w3433_v;
	wire v_w970_v;
	wire v_w5204_v;
	wire v_w4573_v;
	wire v_w6156_v;
	wire v_w1463_v;
	wire v_w5766_v;
	wire v_w2202_v;
	wire v_w7868_v;
	wire v_w7712_v;
	wire v_w1854_v;
	wire v_w3077_v;
	wire v_w6698_v;
	wire v_w737_v;
	wire v_w7903_v;
	wire v_w2755_v;
	wire v_w3147_v;
	wire v_w2155_v;
	wire v_w5798_v;
	wire v_w967_v;
	wire v_w2337_v;
	wire v_w7502_v;
	wire v_w6626_v;
	wire v_w7573_v;
	wire v_w7666_v;
	wire v_w2827_v;
	wire v_w7095_v;
	wire v_w699_v;
	wire v_w2675_v;
	wire v_w4295_v;
	wire v_w409_v;
	wire v_w2073_v;
	wire v_w4199_v;
	reg v_s72_v;
	wire v_w2951_v;
	wire v_w7_v;
	wire v_w2811_v;
	wire v_w209_v;
	wire v_w7322_v;
	wire v_w5064_v;
	wire v_w4886_v;
	wire v_w4826_v;
	wire v_w7155_v;
	wire v_w4164_v;
	wire v_w5783_v;
	wire v_w3334_v;
	wire v_w5125_v;
	wire v_w5933_v;
	wire v_w3471_v;
	wire v_w4511_v;
	wire v_w7973_v;
	wire v_w4601_v;
	wire v_w3652_v;
	wire v_w381_v;
	wire v_w6351_v;
	wire v_w2742_v;
	wire v_w2359_v;
	wire v_w382_v;
	wire v_w4591_v;
	wire v_w6518_v;
	wire v_w886_v;
	wire v_w2149_v;
	wire v_w5287_v;
	wire v_w2434_v;
	wire v_w6059_v;
	wire v_w2550_v;
	wire v_w6566_v;
	wire v_w6295_v;
	wire v_w5072_v;
	wire v_w2612_v;
	wire v_w4366_v;
	wire v_w6539_v;
	wire v_w2946_v;
	wire v_w3037_v;
	wire v_w232_v;
	wire v_w8251_v;
	wire v_w5284_v;
	wire v_w254_v;
	reg v_s495_v;
	wire v_w6781_v;
	wire v_w3528_v;
	wire v_w178_v;
	wire v_w3702_v;
	wire v_w936_v;
	wire v_w3646_v;
	wire v_w6723_v;
	wire v_w4378_v;
	reg v_s222_v;
	wire v_w6585_v;
	wire v_w7016_v;
	wire v_w2547_v;
	wire v_w163_v;
	wire v_w2223_v;
	wire v_w139_v;
	reg v_s79_v;
	reg v_s247_v;
	reg v_s472_v;
	wire v_w6036_v;
	wire v_w6113_v;
	wire v_w21_v;
	wire v_w7687_v;
	wire v_w7749_v;
	wire v_w5212_v;
	wire v_w4213_v;
	wire v_w2227_v;
	wire v_w884_v;
	wire v_w1749_v;
	wire v_w784_v;
	wire v_w6342_v;
	wire v_w7185_v;
	wire v_w6930_v;
	wire v_w7619_v;
	wire v_w1713_v;
	wire v_w488_v;
	wire v_w7959_v;
	wire v_w4763_v;
	wire v_w7221_v;
	wire v_w4953_v;
	wire v_w663_v;
	wire v_w2895_v;
	wire v_w1222_v;
	wire v_w7995_v;
	wire v_w2848_v;
	wire v_w5047_v;
	wire v_w152_v;
	wire v_w806_v;
	wire v_w1151_v;
	wire v_w7980_v;
	wire v_w1332_v;
	wire v_w3301_v;
	wire v_w4609_v;
	wire v_w7286_v;
	wire v_w6476_v;
	reg v_s487_v;
	wire v_w283_v;
	wire v_w2454_v;
	wire v_w7998_v;
	wire v_w5815_v;
	wire v_w4845_v;
	wire v_w4906_v;
	wire v_w7691_v;
	wire v_w1089_v;
	wire v_w3216_v;
	wire v_w1946_v;
	wire v_w817_v;
	wire v_w149_v;
	wire v_w105_v;
	wire v_w3908_v;
	wire v_w1300_v;
	wire v_w1675_v;
	wire v_w7700_v;
	wire v_w7692_v;
	wire v_w2923_v;
	wire v_w4303_v;
	wire v_w4944_v;
	wire v_w3995_v;
	wire v_w5376_v;
	wire v_w474_v;
	wire v_w869_v;
	wire v_w4765_v;
	wire v_w6180_v;
	wire v_w556_v;
	wire v_w8157_v;
	wire v_w7856_v;
	wire v_w6889_v;
	wire v_w5684_v;
	wire v_w4777_v;
	wire v_w1993_v;
	wire v_w2889_v;
	wire v_w6804_v;
	wire v_w293_v;
	reg v_s435_v;
	wire v_w4519_v;
	wire v_w5958_v;
	wire v_w6122_v;
	wire v_w3823_v;
	wire v_w5398_v;
	reg v_s394_v;
	wire v_w5908_v;
	wire v_w2086_v;
	wire v_w43_v;
	wire v_w2653_v;
	wire v_w685_v;
	wire v_w4040_v;
	wire v_w6097_v;
	wire v_w6937_v;
	wire v_w3848_v;
	wire v_w7066_v;
	wire v_w8000_v;
	wire v_w7015_v;
	wire v_w2575_v;
	reg v_s287_v;
	wire v_w7595_v;
	wire v_w4856_v;
	wire v_w984_v;
	wire v_w7547_v;
	wire v_w3295_v;
	wire v_w415_v;
	wire v_w2257_v;
	wire v_w4459_v;
	wire v_w4398_v;
	wire v_w4718_v;
	wire v_w4059_v;
	wire v_w3222_v;
	reg v_s31_v;
	wire v_w7432_v;
	wire v_w5258_v;
	reg v_s457_v;
	wire v_w5942_v;
	wire v_w5448_v;
	wire v_w520_v;
	wire v_w2404_v;
	wire v_w1326_v;
	reg v_s271_v;
	wire v_w1886_v;
	wire v_w3184_v;
	wire v_w2117_v;
	wire v_w2077_v;
	wire v_w3005_v;
	wire v_w4222_v;
	wire v_w173_v;
	wire v_w687_v;
	wire v_w2196_v;
	wire v_w3838_v;
	wire v_w2733_v;
	wire v_w3797_v;
	wire v_w7624_v;
	wire v_w5493_v;
	reg v_s158_v;
	wire v_w3755_v;
	wire v_w271_v;
	wire v_w4457_v;
	wire v_w1207_v;
	wire v_w3451_v;
	wire v_w6578_v;
	wire v_w4654_v;
	wire v_w3950_v;
	wire v_w3127_v;
	wire v_w6760_v;
	wire v_w4318_v;
	wire v_w2071_v;
	wire v_w7279_v;
	wire v_w6021_v;
	wire v_w1251_v;
	reg v_s241_v;
	wire v_w5438_v;
	wire v_w6556_v;
	wire v_w6699_v;
	wire v_w4895_v;
	wire v_w3225_v;
	reg v_s61_v;
	wire v_w7618_v;
	wire v_w7782_v;
	wire v_w5653_v;
	wire v_w3057_v;
	wire v_w4513_v;
	reg v_s492_v;
	wire v_w4966_v;
	wire v_w192_v;
	wire v_w3220_v;
	wire v_w1798_v;
	wire v_w5621_v;
	wire v_w4780_v;
	wire v_w3042_v;
	wire v_w920_v;
	wire v_w1965_v;
	wire v_w4540_v;
	wire v_w5616_v;
	wire v_w5230_v;
	wire v_w270_v;
	wire v_w5465_v;
	wire v_w5651_v;
	wire v_w1778_v;
	wire v_w5089_v;
	wire v_w7512_v;
	wire v_w2458_v;
	wire v_w2524_v;
	wire v_w620_v;
	wire v_w211_v;
	wire v_w3798_v;
	wire v_w2064_v;
	wire v_w388_v;
	wire v_w4325_v;
	wire v_w3895_v;
	wire v_w1446_v;
	wire v_w2959_v;
	wire v_w6086_v;
	wire v_w4104_v;
	wire v_w4629_v;
	wire v_w8085_v;
	wire v_w4030_v;
	wire v_w4604_v;
	wire v_w7574_v;
	wire v_w162_v;
	wire v_w7896_v;
	reg v_s184_v;
	wire v_w2769_v;
	wire v_w5710_v;
	wire v_w6244_v;
	wire v_w1751_v;
	wire v_w4727_v;
	wire v_w5927_v;
	wire v_w3281_v;
	wire v_w7872_v;
	wire v_w4255_v;
	wire v_w7104_v;
	wire v_o15_v;
	wire v_w5559_v;
	wire v_w7217_v;
	wire v_w1964_v;
	wire v_w1911_v;
	wire v_w4761_v;
	wire v_w7966_v;
	wire v_w7267_v;
	wire v_w2111_v;
	wire v_w276_v;
	wire v_w3571_v;
	wire v_w3930_v;
	wire v_w3272_v;
	wire v_w5601_v;
	wire v_w1454_v;
	wire v_w824_v;
	wire v_w3169_v;
	wire v_w2904_v;
	wire v_w2025_v;
	wire v_w4241_v;
	wire v_w7142_v;
	wire v_w7197_v;
	wire v_w4026_v;
	wire v_w969_v;
	wire v_w4484_v;
	wire v_w7077_v;
	wire v_w3573_v;
	wire v_w3751_v;
	wire v_w1819_v;
	wire v_w842_v;
	reg v_s368_v;
	wire v_w2157_v;
	wire v_w6329_v;
	wire v_w1608_v;
	wire v_w811_v;
	wire v_w5711_v;
	wire v_w4052_v;
	wire v_w1830_v;
	wire v_w2104_v;
	wire v_w4887_v;
	wire v_w7330_v;
	wire v_w8224_v;
	wire v_w58_v;
	wire v_w517_v;
	wire v_w2795_v;
	wire v_w333_v;
	wire v_w6709_v;
	wire v_w5536_v;
	wire v_w5246_v;
	reg v_s490_v;
	wire v_w7552_v;
	wire v_w2844_v;
	wire v_w8083_v;
	wire v_w6783_v;
	wire v_w1844_v;
	wire v_w2123_v;
	wire v_w2913_v;
	wire v_w2396_v;
	wire v_w1283_v;
	wire v_w7950_v;
	wire v_w7779_v;
	wire v_w6365_v;
	wire v_w7912_v;
	wire v_w2098_v;
	wire v_w2116_v;
	wire v_w5346_v;
	wire v_w7161_v;
	wire v_w4536_v;
	wire v_w700_v;
	wire v_w6913_v;
	wire v_w593_v;
	wire v_w1490_v;
	wire v_w5596_v;
	wire v_w1256_v;
	wire v_w505_v;
	wire v_w5005_v;
	wire v_w4031_v;
	wire v_w2105_v;
	wire v_w6643_v;
	wire v_w1590_v;
	wire v_w7586_v;
	wire v_w6044_v;
	wire v_w3458_v;
	wire v_w4188_v;
	wire v_w7770_v;
	wire v_w1926_v;
	wire v_w4427_v;
	wire v_w7873_v;
	wire v_w3231_v;
	reg v_s7_v;
	wire v_w2563_v;
	wire v_w458_v;
	wire v_w3942_v;
	wire v_w7018_v;
	wire v_w622_v;
	wire v_w7521_v;
	wire v_w5009_v;
	wire v_w8180_v;
	wire v_w7461_v;
	wire v_w4203_v;
	wire v_w1670_v;
	wire v_w1096_v;
	wire v_w904_v;
	wire v_w56_v;
	wire v_w4998_v;
	wire v_w8232_v;
	reg v_s208_v;
	wire v_w2681_v;
	wire v_w2474_v;
	wire v_w2830_v;
	wire v_w5114_v;
	reg v_s106_v;
	wire v_w3637_v;
	wire v_w598_v;
	wire v_w4259_v;
	wire v_w5788_v;
	wire v_w3974_v;
	wire v_w4667_v;
	wire v_w1905_v;
	wire v_w1059_v;
	wire v_w4339_v;
	wire v_w5341_v;
	wire v_w5315_v;
	wire v_w7925_v;
	wire v_w696_v;
	wire v_w8048_v;
	wire v_w2328_v;
	wire v_w1609_v;
	wire v_w4206_v;
	wire v_w4608_v;
	wire v_w3261_v;
	reg v_s14_v;
	wire v_w5173_v;
	wire v_w434_v;
	wire v_w4082_v;
	wire v_w5606_v;
	wire v_w6359_v;
	wire v_w5403_v;
	wire v_w2409_v;
	wire v_w6383_v;
	wire v_w7009_v;
	wire v_w1790_v;
	wire v_w3499_v;
	wire v_w6075_v;
	wire v_w6998_v;
	wire v_w3828_v;
	wire v_w8065_v;
	wire v_w8138_v;
	wire v_w4210_v;
	wire v_w5907_v;
	wire v_w1377_v;
	wire v_w7041_v;
	wire v_w1999_v;
	wire v_w703_v;
	wire v_w3257_v;
	wire v_w6163_v;
	wire v_w5062_v;
	wire v_w4179_v;
	wire v_w5317_v;
	wire v_w3123_v;
	wire v_w4069_v;
	wire v_w823_v;
	wire v_w5795_v;
	wire v_w5929_v;
	wire v_w1217_v;
	wire v_w6270_v;
	wire v_w5898_v;
	wire v_w4218_v;
	wire v_w137_v;
	wire v_w6784_v;
	wire v_w3101_v;
	wire v_w5625_v;
	reg v_s399_v;
	wire v_w6202_v;
	reg v_s507_v;
	wire v_w133_v;
	wire v_w1616_v;
	wire v_w603_v;
	wire v_w4352_v;
	wire v_w2399_v;
	wire v_w7919_v;
	wire v_w5899_v;
	wire v_w3322_v;
	wire v_w88_v;
	wire v_w7611_v;
	wire v_w4006_v;
	wire v_w2150_v;
	wire v_w431_v;
	wire v_w4346_v;
	wire v_w4595_v;
	reg v_s420_v;
	wire v_w2760_v;
	wire v_w6080_v;
	wire v_w6667_v;
	wire v_w5610_v;
	wire v_w7118_v;
	wire v_w2500_v;
	wire v_w7813_v;
	wire v_w1320_v;
	wire v_w625_v;
	wire v_w1606_v;
	wire v_w816_v;
	wire v_w6927_v;
	wire v_w1991_v;
	wire v_w4681_v;
	wire v_w3389_v;
	reg v_s141_v;
	wire v_w369_v;
	wire v_w1427_v;
	wire v_w1178_v;
	wire v_w5466_v;
	wire v_w4957_v;
	wire v_w2762_v;
	wire v_w2692_v;
	wire v_w4343_v;
	wire v_w1657_v;
	wire v_w3485_v;
	wire v_w1040_v;
	wire v_w8141_v;
	wire v_w348_v;
	wire v_w3382_v;
	wire v_w2767_v;
	wire v_w1142_v;
	wire v_w127_v;
	wire v_w309_v;
	wire v_w7058_v;
	wire v_w375_v;
	wire v_w4864_v;
	wire v_w6926_v;
	wire v_w7403_v;
	wire v_w4790_v;
	wire v_w6239_v;
	wire v_w1508_v;
	wire v_w2996_v;
	wire v_w4521_v;
	wire v_w6490_v;
	wire v_w3683_v;
	wire v_w6146_v;
	wire v_w326_v;
	wire v_w4492_v;
	wire v_w228_v;
	wire v_w7311_v;
	wire v_w7549_v;
	wire v_w4420_v;
	wire v_w6407_v;
	wire v_w310_v;
	wire v_w7121_v;
	wire v_w6911_v;
	wire v_w5074_v;
	wire v_w6632_v;
	wire v_w6618_v;
	wire v_w944_v;
	wire v_w3251_v;
	wire v_w2604_v;
	wire v_w2118_v;
	wire v_w4881_v;
	reg v_s259_v;
	wire v_w988_v;
	wire v_w1381_v;
	wire v_w4798_v;
	wire v_w5443_v;
	wire v_w3682_v;
	wire v_w5537_v;
	wire v_w7034_v;
	wire v_w6052_v;
	wire v_w4025_v;
	wire v_w6233_v;
	wire v_w3714_v;
	wire v_w6928_v;
	wire v_w6931_v;
	wire v_w7953_v;
	wire v_w7294_v;
	wire v_w5737_v;
	wire v_w6521_v;
	wire v_w5412_v;
	wire v_w5104_v;
	wire v_w8131_v;
	wire v_w1692_v;
	wire v_w1862_v;
	wire v_w4830_v;
	wire v_w3981_v;
	wire v_w2302_v;
	wire v_w1931_v;
	wire v_w7135_v;
	wire v_w7316_v;
	wire v_w2315_v;
	wire v_w3287_v;
	wire v_w4436_v;
	wire v_w7808_v;
	wire v_w5880_v;
	wire v_w2813_v;
	wire v_w3698_v;
	wire v_w7888_v;
	wire v_w4347_v;
	reg v_s23_v;
	wire v_w1246_v;
	wire v_w6609_v;
	wire v_w4551_v;
	wire v_w3338_v;
	wire v_w3665_v;
	wire v_w5564_v;
	wire v_w6983_v;
	wire v_w5440_v;
	reg v_s104_v;
	wire v_w2087_v;
	wire v_w6330_v;
	wire v_w765_v;
	wire v_w923_v;
	wire v_w7177_v;
	wire v_w3706_v;
	wire v_w2175_v;
	wire v_w6509_v;
	wire v_w4768_v;
	wire v_w1227_v;
	wire v_w5053_v;
	wire v_w3678_v;
	wire v_w159_v;
	wire v_w7093_v;
	reg v_s248_v;
	wire v_w1643_v;
	wire v_w217_v;
	wire v_w6218_v;
	wire v_w7275_v;
	reg v_s246_v;
	wire v_w3487_v;
	reg v_s69_v;
	wire v_w7858_v;
	wire v_w6831_v;
	wire v_w3391_v;
	reg v_s503_v;
	wire v_w2716_v;
	wire v_w6403_v;
	wire v_w5759_v;
	wire v_w5518_v;
	wire v_w2747_v;
	wire v_w3358_v;
	wire v_w7506_v;
	wire v_w5121_v;
	wire v_w2016_v;
	wire v_w6812_v;
	wire v_w5800_v;
	wire v_w8005_v;
	wire v_w606_v;
	wire v_w5966_v;
	wire v_w1415_v;
	wire v_w5260_v;
	wire v_w5889_v;
	wire v_w2156_v;
	wire v_w4442_v;
	wire v_w1273_v;
	wire v_w3080_v;
	reg v_s265_v;
	wire v_w4501_v;
	wire v_w7793_v;
	wire v_w6640_v;
	wire v_w7891_v;
	wire v_w3277_v;
	wire v_w952_v;
	wire v_w2381_v;
	wire v_w4399_v;
	wire v_w6891_v;
	wire v_w4284_v;
	wire v_w6223_v;
	wire v_w3633_v;
	wire v_w7865_v;
	wire v_w2414_v;
	wire v_w5887_v;
	reg v_s286_v;
	wire v_w1553_v;
	wire v_w4739_v;
	wire v_w3636_v;
	wire v_w7939_v;
	wire v_w5374_v;
	wire v_w1367_v;
	wire v_w6285_v;
	wire v_w7659_v;
	wire v_w2643_v;
	wire v_w3130_v;
	wire v_w7368_v;
	wire v_w4842_v;
	wire v_w6249_v;
	wire v_w2866_v;
	wire v_w2437_v;
	wire v_w7927_v;
	wire v_w7800_v;
	wire v_w8024_v;
	wire v_w2052_v;
	wire v_w5857_v;
	wire v_w3079_v;
	wire v_w4938_v;
	wire v_w971_v;
	wire v_w2037_v;
	wire v_w3454_v;
	wire v_w8150_v;
	wire v_w3687_v;
	wire v_w8201_v;
	reg v_s258_v;
	wire v_w1593_v;
	wire v_w8118_v;
	wire v_w6184_v;
	wire v_w4070_v;
	wire v_w5558_v;
	wire v_w1144_v;
	wire v_w6906_v;
	wire v_w4602_v;
	wire v_w7735_v;
	wire v_w7249_v;
	wire v_w6363_v;
	wire v_w6390_v;
	wire v_w615_v;
	wire v_w4289_v;
	wire v_w7943_v;
	wire v_w7748_v;
	wire v_w480_v;
	wire v_w7012_v;
	reg v_s253_v;
	wire v_w1189_v;
	wire v_w2939_v;
	wire v_w710_v;
	wire v_w4542_v;
	wire v_w734_v;
	wire v_w7083_v;
	wire v_w7592_v;
	wire v_w8115_v;
	wire v_w5020_v;
	wire v_w8165_v;
	wire v_w7054_v;
	wire v_w3245_v;
	wire v_w1705_v;
	wire v_w5560_v;
	wire v_w2859_v;
	wire v_w7725_v;
	wire v_w29_v;
	wire v_w2332_v;
	wire v_w5357_v;
	wire v_w8155_v;
	wire v_w6530_v;
	wire v_w2254_v;
	wire v_w4499_v;
	wire v_w1465_v;
	wire v_w3342_v;
	wire v_w7850_v;
	wire v_w2717_v;
	wire v_w3045_v;
	wire v_w5078_v;
	wire v_w3076_v;
	wire v_w6557_v;
	wire v_w2400_v;
	wire v_w6701_v;
	wire v_w3016_v;
	wire v_w8214_v;
	wire v_w6131_v;
	wire v_w4105_v;
	wire v_w3590_v;
	wire v_w3297_v;
	wire v_w6642_v;
	wire v_w4972_v;
	wire v_w5268_v;
	wire v_w658_v;
	wire v_w2229_v;
	wire v_w4435_v;
	wire v_w2503_v;
	wire v_w439_v;
	wire v_w2932_v;
	wire v_w4429_v;
	wire v_w4925_v;
	reg v_s389_v;
	wire v_w2240_v;
	wire v_w4432_v;
	wire v_w3614_v;
	wire v_w6670_v;
	wire v_w2857_v;
	wire v_w4580_v;
	wire v_w4933_v;
	wire v_w6398_v;
	wire v_w1047_v;
	wire v_w2689_v;
	wire v_w7660_v;
	wire v_w7241_v;
	wire v_w7179_v;
	wire v_w6307_v;
	wire v_w1554_v;
	wire v_w7964_v;
	wire v_w4899_v;
	wire v_w626_v;
	wire v_w4410_v;
	wire v_w1061_v;
	wire v_w5257_v;
	wire v_w535_v;
	wire v_w3365_v;
	wire v_w7920_v;
	wire v_w142_v;
	wire v_w7303_v;
	wire v_w2888_v;
	wire v_w6198_v;
	wire v_w2394_v;
	wire v_w363_v;
	wire v_w4841_v;
	wire v_w1493_v;
	wire v_w5026_v;
	wire v_w493_v;
	wire v_w4455_v;
	wire v_w1866_v;
	wire v_w1472_v;
	reg v_s266_v;
	reg v_s77_v;
	wire v_w6715_v;
	wire v_w5065_v;
	wire v_w3210_v;
	wire v_w1591_v;
	wire v_w3400_v;
	wire v_w531_v;
	reg v_s64_v;
	wire v_w829_v;
	wire v_w536_v;
	wire v_w3512_v;
	wire v_w4840_v;
	wire v_w3001_v;
	wire v_w808_v;
	wire v_w1681_v;
	wire v_w7056_v;
	wire v_w5691_v;
	wire v_w2539_v;
	reg v_s80_v;
	wire v_w3812_v;
	wire v_w2329_v;
	wire v_w6090_v;
	wire v_w6547_v;
	wire v_w1045_v;
	wire v_w2024_v;
	wire v_w5840_v;
	wire v_w299_v;
	wire v_w3519_v;
	wire v_w3649_v;
	wire v_w4317_v;
	wire v_w2447_v;
	wire v_w6322_v;
	wire v_w8110_v;
	wire v_w411_v;
	wire v_w6858_v;
	wire v_w762_v;
	wire v_w2049_v;
	wire v_w2933_v;
	wire v_w7216_v;
	reg v_s237_v;
	wire v_w3996_v;
	wire v_w2208_v;
	wire v_w3332_v;
	wire v_w4228_v;
	wire v_w5973_v;
	reg v_s68_v;
	reg v_s341_v;
	wire v_w3348_v;
	wire v_w3428_v;
	wire v_w7754_v;
	wire v_w2059_v;
	wire v_w144_v;
	wire v_w3885_v;
	wire v_w8_v;
	wire v_w756_v;
	wire v_w6177_v;
	wire v_w7116_v;
	wire v_w5514_v;
	wire v_w2010_v;
	wire v_w2704_v;
	wire v_w1318_v;
	wire v_w1555_v;
	wire v_w5924_v;
	reg v_s500_v;
	wire v_w402_v;
	wire v_w5250_v;
	wire v_w6037_v;
	wire v_w6119_v;
	wire v_w2100_v;
	wire v_w2581_v;
	wire v_w5793_v;
	reg v_s363_v;
	wire v_w6427_v;
	wire v_w1462_v;
	reg v_s440_v;
	wire v_w7665_v;
	wire v_w5154_v;
	wire v_w4593_v;
	wire v_w1310_v;
	wire v_w5743_v;
	reg v_s313_v;
	wire v_w3031_v;
	wire v_w5479_v;
	wire v_w5728_v;
	wire v_w2242_v;
	wire v_w805_v;
	wire v_w3530_v;
	wire v_w5916_v;
	wire v_w6039_v;
	wire v_w1641_v;
	wire v_w7188_v;
	wire v_w931_v;
	wire v_w7489_v;
	wire v_w5789_v;
	wire v_w8034_v;
	wire v_w5411_v;
	wire v_w3656_v;
	wire v_w3349_v;
	wire v_w3183_v;
	wire v_w4143_v;
	wire v_w4943_v;
	wire v_w6755_v;
	wire v_w3928_v;
	wire v_w6997_v;
	wire v_w1402_v;
	wire v_w856_v;
	wire v_w7658_v;
	wire v_w5843_v;
	wire v_w4426_v;
	reg v_s109_v;
	wire v_w7822_v;
	wire v_w374_v;
	wire v_w6933_v;
	wire v_w242_v;
	wire v_w4858_v;
	wire v_w5431_v;
	wire v_w713_v;
	reg v_s34_v;
	wire v_w4639_v;
	wire v_w5579_v;
	wire v_w5458_v;
	wire v_w4583_v;
	wire v_w1438_v;
	wire v_w6854_v;
	wire v_w1536_v;
	wire v_w3630_v;
	wire v_w1780_v;
	wire v_w366_v;
	wire v_w3911_v;
	reg v_s342_v;
	wire v_w4365_v;
	wire v_w6975_v;
	wire v_w5782_v;
	wire v_w4940_v;
	wire v_w264_v;
	wire v_w5067_v;
	wire v_w2910_v;
	wire v_w2363_v;
	wire v_w7823_v;
	wire v_w2702_v;
	wire v_w3566_v;
	wire v_w5854_v;
	wire v_w7419_v;
	wire v_w5890_v;
	reg v_s403_v;
	wire v_w4852_v;
	wire v_w3346_v;
	wire v_w2478_v;
	wire v_w3926_v;
	wire v_w1956_v;
	wire v_w2960_v;
	wire v_w3833_v;
	wire v_w7738_v;
	wire v_w8095_v;
	wire v_w4445_v;
	wire v_w6291_v;
	wire v_w3923_v;
	wire v_w7883_v;
	wire v_w7609_v;
	wire v_w601_v;
	wire v_w4139_v;
	wire v_w6101_v;
	wire v_w3011_v;
	wire v_w4816_v;
	wire v_w4482_v;
	wire v_w7346_v;
	wire v_w3874_v;
	wire v_w7932_v;
	wire v_w7490_v;
	wire v_w868_v;
	wire v_w6679_v;
	reg v_s96_v;
	wire v_w3237_v;
	wire v_w3097_v;
	wire v_w7205_v;
	wire v_w7392_v;
	wire v_w7430_v;
	wire v_w2849_v;
	wire v_w5813_v;
	wire v_w1560_v;
	wire v_w1729_v;
	wire v_w6912_v;
	wire v_w6850_v;
	wire v_w1777_v;
	wire v_w7484_v;
	wire v_w7528_v;
	wire v_w6002_v;
	wire v_w2679_v;
	wire v_w1066_v;
	wire v_w3199_v;
	wire v_w4390_v;
	reg v_s199_v;
	wire v_w837_v;
	wire v_w3276_v;
	wire v_w5523_v;
	wire v_w5632_v;
	wire v_w7295_v;
	wire v_w2085_v;
	wire v_w504_v;
	wire v_w8200_v;
	wire v_w796_v;
	wire v_w399_v;
	wire v_w2892_v;
	wire v_w4407_v;
	wire v_w5167_v;
	wire v_w7933_v;
	wire v_w128_v;
	wire v_w8098_v;
	wire v_w8047_v;
	wire v_w6697_v;
	wire v_w950_v;
	wire v_w5456_v;
	wire v_w19_v;
	wire v_w6901_v;
	wire v_w3871_v;
	wire v_w6338_v;
	reg v_s118_v;
	wire v_w84_v;
	wire v_w1416_v;
	wire v_w5644_v;
	wire v_w2426_v;
	wire v_w2193_v;
	wire v_w1686_v;
	wire v_w913_v;
	wire v_w7397_v;
	wire v_w15_v;
	wire v_w1934_v;
	wire v_w629_v;
	wire v_w6414_v;
	reg v_s274_v;
	wire v_w7817_v;
	wire v_w2408_v;
	reg v_s226_v;
	wire v_w5303_v;
	wire v_w1791_v;
	wire v_w3296_v;
	wire v_w1788_v;
	reg v_s82_v;
	wire v_w6148_v;
	wire v_w1963_v;
	wire v_w3865_v;
	wire v_w1871_v;
	wire v_w925_v;
	wire v_w2313_v;
	wire v_w7636_v;
	wire v_w1588_v;
	wire v_w8239_v;
	wire v_w6676_v;
	wire v_w4223_v;
	wire v_w184_v;
	wire v_w421_v;
	wire v_w3056_v;
	wire v_w1041_v;
	wire v_w8062_v;
	wire v_w2903_v;
	wire v_w5989_v;
	wire v_w3262_v;
	wire v_w1661_v;
	wire v_w3360_v;
	wire v_w3658_v;
	reg v_s458_v;
	wire v_w8196_v;
	wire v_w3907_v;
	wire v_w7620_v;
	wire v_w5390_v;
	wire v_w250_v;
	wire v_w3260_v;
	wire v_w6834_v;
	wire v_w405_v;
	wire v_w5998_v;
	wire v_w3213_v;
	wire v_w3386_v;
	wire v_w7415_v;
	wire v_w6855_v;
	wire v_w4024_v;
	wire v_w5328_v;
	wire v_w5055_v;
	wire v_w8225_v;
	wire v_o17_v;
	wire v_w4945_v;
	wire v_w4448_v;
	reg v_s279_v;
	wire v_w960_v;
	wire v_w5015_v;
	wire v_w3221_v;
	wire v_w7105_v;
	wire v_w5051_v;
	wire v_w6115_v;
	wire v_w2122_v;
	wire v_w2522_v;
	wire v_w24_v;
	wire v_w8198_v;
	wire v_w5446_v;
	wire v_w4770_v;
	wire v_w342_v;
	wire v_w5694_v;
	wire v_w7094_v;
	wire v_w1159_v;
	wire v_w2828_v;
	wire v_w8011_v;
	wire v_w8145_v;
	wire v_w1226_v;
	wire v_w3164_v;
	wire v_w7762_v;
	wire v_w3388_v;
	wire v_w4592_v;
	wire v_w5439_v;
	wire v_w393_v;
	wire v_w6789_v;
	wire v_w571_v;
	wire v_w3767_v;
	wire v_w1610_v;
	wire v_w5198_v;
	wire v_w4_v;
	wire v_w3052_v;
	wire v_w7644_v;
	wire v_w3477_v;
	wire v_w4391_v;
	wire v_w5723_v;
	wire v_w6500_v;
	wire v_w7013_v;
	wire v_w1435_v;
	wire v_w161_v;
	wire v_w5308_v;
	wire v_w4648_v;
	wire v_w5715_v;
	wire v_w7690_v;
	wire v_w2881_v;
	wire v_w7763_v;
	wire v_w1863_v;
	wire v_w7373_v;
	wire v_w7442_v;
	wire v_w1954_v;
	wire v_w125_v;
	wire v_w5132_v;
	wire v_w3243_v;
	wire v_w870_v;
	wire v_w2845_v;
	reg v_s423_v;
	wire v_w7737_v;
	wire v_w1923_v;
	wire v_w203_v;
	wire v_w3734_v;
	wire v_w65_v;
	wire v_w7000_v;
	wire v_w1386_v;
	reg v_s491_v;
	wire v_w5879_v;
	wire v_w3916_v;
	wire v_w2326_v;
	wire v_w1302_v;
	wire v_w5920_v;
	wire v_w3022_v;
	wire v_w6166_v;
	wire v_w6003_v;
	wire v_w2737_v;
	wire v_w2798_v;
	wire v_w3518_v;
	wire v_w2846_v;
	wire v_w2669_v;
	wire v_w7224_v;
	wire v_w1_v;
	wire v_w5207_v;
	wire v_w2552_v;
	wire v_w6380_v;
	wire v_w2035_v;
	wire v_w993_v;
	wire v_w3207_v;
	reg v_s186_v;
	wire v_w5013_v;
	reg v_s38_v;
	wire v_w6457_v;
	wire v_w5302_v;
	wire v_w1442_v;
	wire v_w6255_v;
	reg v_s240_v;
	wire v_w5462_v;
	wire v_w1138_v;
	wire v_w1764_v;
	wire v_w850_v;
	wire v_w5060_v;
	wire v_w2850_v;
	wire v_w3657_v;
	wire v_w3948_v;
	wire v_w4171_v;
	wire v_w398_v;
	wire v_w2266_v;
	wire v_w2885_v;
	wire v_w1543_v;
	wire v_w4716_v;
	wire v_w3965_v;
	wire v_w2430_v;
	wire v_w4161_v;
	wire v_w351_v;
	wire v_w5007_v;
	wire v_w6974_v;
	wire v_w8192_v;
	wire v_w7138_v;
	wire v_w2192_v;
	wire v_w5846_v;
	wire v_w7518_v;
	wire v_w2_v;
	wire v_w182_v;
	wire v_w4996_v;
	reg v_s257_v;
	wire v_w5295_v;
	wire v_w5050_v;
	wire v_w2564_v;
	reg v_s356_v;
	wire v_w5816_v;
	wire v_w4175_v;
	wire v_w5935_v;
	wire v_w1917_v;
	wire v_w2724_v;
	wire v_w4375_v;
	wire v_w2854_v;
	wire v_w36_v;
	wire v_w977_v;
	wire v_w7365_v;
	wire v_w4282_v;
	wire v_w8076_v;
	wire v_w3770_v;
	wire v_w8170_v;
	wire v_w5981_v;
	wire v_w6658_v;
	wire v_w5987_v;
	wire v_w3606_v;
	reg v_s520_v;
	wire v_w5868_v;
	wire v_w2379_v;
	wire v_w1039_v;
	wire v_w5874_v;
	wire v_w6062_v;
	wire v_w3196_v;
	wire v_w274_v;
	wire v_w1168_v;
	reg v_s484_v;
	wire v_w6396_v;
	wire v_w6675_v;
	wire v_w5228_v;
	wire v_w4611_v;
	wire v_w4876_v;
	wire v_w2520_v;
	wire v_w6717_v;
	wire v_w6835_v;
	wire v_w8166_v;
	wire v_w1716_v;
	wire v_w5735_v;
	reg v_s107_v;
	wire v_w6128_v;
	wire v_w422_v;
	wire v_w7947_v;
	wire v_w7398_v;
	wire v_w645_v;
	wire v_w5797_v;
	wire v_w6773_v;
	wire v_w5340_v;
	wire v_w2940_v;
	wire v_w2576_v;
	wire v_w650_v;
	wire v_w7520_v;
	wire v_w7811_v;
	wire v_w8119_v;
	wire v_w5116_v;
	wire v_w2636_v;
	wire v_w2816_v;
	wire v_w9_v;
	wire v_w3548_v;
	wire v_w560_v;
	reg v_s307_v;
	wire v_w5094_v;
	wire v_w3533_v;
	wire v_w5799_v;
	wire v_w1537_v;
	reg v_s187_v;
	wire v_w2551_v;
	wire v_w5354_v;
	wire v_w3364_v;
	wire v_w2219_v;
	reg v_s483_v;
	wire v_w7557_v;
	wire v_w7962_v;
	wire v_w7803_v;
	wire v_w1193_v;
	wire v_w6662_v;
	wire v_w8007_v;
	wire v_w482_v;
	wire v_w2984_v;
	wire v_w1627_v;
	wire v_w4814_v;
	wire v_w2044_v;
	wire v_w5827_v;
	wire v_w2825_v;
	wire v_w4968_v;
	wire v_w6579_v;
	reg v_s366_v;
	wire v_w4081_v;
	wire v_w6412_v;
	wire v_w2967_v;
	wire v_w7204_v;
	wire v_w3553_v;
	wire v_w2560_v;
	wire v_w1779_v;
	wire v_w6767_v;
	wire v_w2457_v;
	wire v_w4148_v;
	wire v_w6512_v;
	wire v_w272_v;
	reg v_s448_v;
	reg v_s192_v;
	wire v_w4470_v;
	wire v_w7560_v;
	wire v_w1071_v;
	wire v_w2046_v;
	wire v_w3643_v;
	wire v_w2648_v;
	wire v_w714_v;
	wire v_w4451_v;
	wire v_w3796_v;
	wire v_w1099_v;
	wire v_w6849_v;
	wire v_w6628_v;
	wire v_w4958_v;
	wire v_w709_v;
	wire v_w2435_v;
	reg v_s209_v;
	wire v_w4607_v;
	wire v_w8030_v;
	wire v_w238_v;
	wire v_w66_v;
	wire v_w5386_v;
	reg v_s362_v;
	wire v_w2917_v;
	wire v_w7526_v;
	wire v_w6159_v;
	wire v_w792_v;
	wire v_w4708_v;
	wire v_w5967_v;
	wire v_w3252_v;
	wire v_w7201_v;
	wire v_w4707_v;
	wire v_w4624_v;
	wire v_w7141_v;
	wire v_w1719_v;
	wire v_w963_v;
	wire v_w6319_v;
	wire v_w7115_v;
	wire v_w3912_v;
	wire v_w1259_v;
	wire v_w2880_v;
	wire v_w4952_v;
	wire v_w451_v;
	wire v_w7694_v;
	wire v_w2777_v;
	wire v_w6644_v;
	wire v_w2405_v;
	wire v_w82_v;
	wire v_w3311_v;
	reg v_s230_v;
	wire v_w1087_v;
	wire v_w2042_v;
	wire v_w4191_v;
	wire v_w2120_v;
	wire v_w741_v;
	reg v_s249_v;
	wire v_w4166_v;
	wire v_w1051_v;
	wire v_w6497_v;
	wire v_w1642_v;
	wire v_w3182_v;
	wire v_w2805_v;
	reg v_s44_v;
	wire v_w6805_v;
	wire v_w6949_v;
	wire v_w6422_v;
	wire v_w6311_v;
	wire v_w3752_v;
	wire v_w6922_v;
	wire v_w6963_v;
	wire v_w3279_v;
	wire v_w3046_v;
	wire v_w4861_v;
	wire v_w4878_v;
	wire v_w775_v;
	wire v_w2255_v;
	wire v_w7167_v;
	wire v_w6206_v;
	wire v_w1784_v;
	wire v_w6287_v;
	wire v_w898_v;
	wire v_w1857_v;
	wire v_w7569_v;
	wire v_w8169_v;
	wire v_w5442_v;
	wire v_w5484_v;
	wire v_w4775_v;
	reg v_s112_v;
	wire v_w5187_v;
	wire v_w3615_v;
	wire v_w1260_v;
	reg v_s89_v;
	wire v_w4817_v;
	wire v_w4075_v;
	wire v_w437_v;
	wire v_w6404_v;
	wire v_w6452_v;
	wire v_w8183_v;
	wire v_w7075_v;
	wire v_w2820_v;
	wire v_w3406_v;
	wire v_w7928_v;
	wire v_w6302_v;
	wire v_w5912_v;
	wire v_w5416_v;
	wire v_w5492_v;
	wire v_w642_v;
	wire v_w3978_v;
	wire v_w707_v;
	wire v_w4898_v;
	wire v_w5659_v;
	wire v_w1908_v;
	wire v_w555_v;
	wire v_w8128_v;
	wire v_w4118_v;
	wire v_w6740_v;
	wire v_w1257_v;
	reg v_s404_v;
	wire v_w5457_v;
	wire v_w6631_v;
	wire v_w5896_v;
	wire v_w8006_v;
	wire v_w5382_v;
	wire v_w6189_v;
	wire v_w3488_v;
	wire v_w8059_v;
	wire v_w8125_v;
	wire v_w4549_v;
	wire v_w7577_v;
	wire v_w6957_v;
	wire v_w3156_v;
	wire v_w4743_v;
	reg v_s262_v;
	wire v_w1601_v;
	wire v_w5732_v;
	wire v_w6645_v;
	wire v_w5436_v;
	wire v_w7073_v;
	wire v_w7313_v;
	wire v_w7632_v;
	wire v_w2937_v;
	wire v_w7570_v;
	wire v_w5613_v;
	wire v_w5451_v;
	wire v_w2148_v;
	wire v_w5818_v;
	wire v_w83_v;
	reg v_s67_v;
	wire v_w1914_v;
	wire v_w5502_v;
	reg v_s468_v;
	wire v_w4802_v;
	wire v_w5294_v;
	wire v_w6173_v;
	wire v_w6323_v;
	wire v_w4752_v;
	wire v_w611_v;
	wire v_w4867_v;
	wire v_w3329_v;
	wire v_w5469_v;
	wire v_w1242_v;
	wire v_w3459_v;
	wire v_w523_v;
	wire v_w2163_v;
	wire v_w1264_v;
	wire v_w5362_v;
	wire v_w6453_v;
	wire v_w1685_v;
	wire v_w3869_v;
	wire v_w3205_v;
	wire v_w3317_v;
	wire v_w1239_v;
	wire v_w4221_v;
	wire v_w6941_v;
	wire v_w2336_v;
	wire v_w3904_v;
	wire v_w2403_v;
	wire v_w2134_v;
	wire v_w2206_v;
	wire v_w1890_v;
	wire v_w6241_v;
	wire v_w6562_v;
	wire v_w7907_v;
	wire v_w5672_v;
	wire v_w5160_v;
	reg v_s111_v;
	wire v_w6260_v;
	wire v_w7832_v;
	wire v_w6235_v;
	wire v_w2456_v;
	wire v_w4096_v;
	wire v_w1299_v;
	wire v_w1707_v;
	wire v_w2555_v;
	wire v_w3762_v;
	wire v_w1483_v;
	wire v_w6099_v;
	wire v_w1747_v;
	wire v_w7348_v;
	reg v_s297_v;
	wire v_w7124_v;
	wire v_w1802_v;
	wire v_w4744_v;
	wire v_w4216_v;
	wire v_w4837_v;
	wire v_w3313_v;
	wire v_w773_v;
	wire v_w3192_v;
	wire v_w5082_v;
	wire v_w1214_v;
	wire v_w6904_v;
	wire v_w2340_v;
	wire v_w4516_v;
	wire v_w3569_v;
	wire v_w3214_v;
	wire v_w4929_v;
	wire v_w3830_v;
	wire v_w3098_v;
	wire v_w1720_v;
	wire v_w6434_v;
	wire v_w7071_v;
	wire v_w5415_v;
	wire v_w6813_v;
	wire v_w5423_v;
	wire v_w3803_v;
	reg v_s424_v;
	wire v_w7369_v;
	wire v_w3899_v;
	wire v_w3891_v;
	wire v_w4638_v;
	wire v_w5805_v;
	wire v_w1653_v;
	reg v_s304_v;
	wire v_w6141_v;
	wire v_w7612_v;
	wire v_w1741_v;
	wire v_w6237_v;
	wire v_w570_v;
	wire v_w6621_v;
	wire v_w3709_v;
	wire v_w3270_v;
	wire v_w4689_v;
	wire v_w2195_v;
	wire v_w3111_v;
	wire v_w1258_v;
	wire v_w6482_v;
	wire v_w6820_v;
	wire v_w976_v;
	wire v_w5130_v;
	wire v_w4960_v;
	wire v_w2958_v;
	wire v_w4281_v;
	wire v_w3527_v;
	wire v_w1987_v;
	wire v_w465_v;
	wire v_w1635_v;
	wire v_w5165_v;
	wire v_w7568_v;
	wire v_w7096_v;
	wire v_w8016_v;
	wire v_w975_v;
	wire v_w4803_v;
	wire v_w3267_v;
	wire v_w3920_v;
	wire v_w487_v;
	wire v_w1107_v;
	wire v_w3310_v;
	wire v_w2860_v;
	wire v_w502_v;
	wire v_w2894_v;
	wire v_w1628_v;
	wire v_w4547_v;
	reg v_s446_v;
	wire v_w1414_v;
	wire v_w6584_v;
	wire v_w5624_v;
	wire v_w3470_v;
	wire v_w3635_v;
	wire v_w1585_v;
	wire v_w8246_v;
	wire v_w1546_v;
	wire v_w5201_v;
	wire v_w294_v;
	wire v_w7198_v;
	wire v_w5676_v;
	wire v_w1431_v;
	wire v_w1126_v;
	wire v_w5546_v;
	wire v_w2966_v;
	wire v_w156_v;
	wire v_w5999_v;
	wire v_w1038_v;
	wire v_w7683_v;
	wire v_w2677_v;
	wire v_w4152_v;
	wire v_w7857_v;
	wire v_w5338_v;
	wire v_w3726_v;
	wire v_w6976_v;
	wire v_w5241_v;
	wire v_w5646_v;
	wire v_w2483_v;
	wire v_w3178_v;
	wire v_w2289_v;
	wire v_w6567_v;
	reg v_s498_v;
	wire v_w5323_v;
	wire v_w793_v;
	wire v_w1838_v;
	wire v_w2479_v;
	wire v_w7605_v;
	wire v_w4786_v;
	wire v_w2189_v;
	wire v_w4149_v;
	reg v_s385_v;
	wire v_w7576_v;
	wire v_w5481_v;
	wire v_w6763_v;
	reg v_s375_v;
	wire v_w6600_v;
	reg v_s62_v;
	wire v_w2053_v;
	wire v_w4340_v;
	wire v_w7827_v;
	wire v_w7225_v;
	wire v_w7450_v;
	wire v_w5604_v;
	wire v_w4610_v;
	wire v_w7308_v;
	wire v_w44_v;
	wire v_w6502_v;
	wire v_w2465_v;
	wire v_w343_v;
	wire v_w2050_v;
	wire v_w7945_v;
	wire v_w651_v;
	wire v_w3574_v;
	wire v_w6592_v;
	wire v_w2654_v;
	wire v_w3244_v;
	wire v_w367_v;
	wire v_w1212_v;
	wire v_w6519_v;
	wire v_w686_v;
	wire v_w2764_v;
	wire v_w6051_v;
	wire v_w5220_v;
	wire v_w1001_v;
	wire v_w2823_v;
	wire v_w3321_v;
	wire v_w5821_v;
	wire v_w8208_v;
	wire v_w5530_v;
	wire v_w7144_v;
	reg v_s331_v;
	wire v_w7603_v;
	wire v_w4538_v;
	wire v_w6892_v;
	wire v_w3480_v;
	wire v_w4425_v;
	wire v_w4275_v;
	reg v_s379_v;
	wire v_w7493_v;
	wire v_w3023_v;
	wire v_w2877_v;
	wire v_w186_v;
	wire v_w4504_v;
	wire v_w6151_v;
	wire v_w563_v;
	wire v_w3860_v;
	wire v_w4581_v;
	wire v_w3559_v;
	wire v_w1978_v;
	wire v_o4_v;
	wire v_w2048_v;
	wire v_w5111_v;
	wire v_w3893_v;
	wire v_w3898_v;
	wire v_w1774_v;
	wire v_w6710_v;
	wire v_w3067_v;
	wire v_w5590_v;
	wire v_w4880_v;
	reg v_s387_v;
	wire v_w2494_v;
	wire v_w5023_v;
	wire v_w6420_v;
	reg v_s438_v;
	wire v_w2542_v;
	wire v_w2342_v;
	wire v_w675_v;
	wire v_w8103_v;
	wire v_w1545_v;
	wire v_w7859_v;
	wire v_w3119_v;
	wire v_w5044_v;
	wire v_w3140_v;
	wire v_w2113_v;
	wire v_w5070_v;
	wire v_w3679_v;
	wire v_w7756_v;
	wire v_w7134_v;
	wire v_w1598_v;
	wire v_w550_v;
	wire v_w6887_v;
	wire v_w2464_v;
	wire v_w2660_v;
	wire v_w7979_v;
	wire v_w527_v;
	wire v_w5093_v;
	wire v_w1953_v;
	wire v_w5043_v;
	wire v_w5831_v;
	wire v_w5944_v;
	wire v_w6480_v;
	wire v_w4351_v;
	wire v_w1042_v;
	wire v_w5222_v;
	wire v_w5807_v;
	wire v_w7425_v;
	wire v_w6350_v;
	wire v_w7523_v;
	wire v_w2354_v;
	wire v_w541_v;
	wire v_w3988_v;
	wire v_w1694_v;
	wire v_w4125_v;
	wire v_w3946_v;
	wire v_w2413_v;
	wire v_w1967_v;
	wire v_w2158_v;
	reg v_s204_v;
	wire v_w7786_v;
	reg v_s508_v;
	wire v_w499_v;
	wire v_w4335_v;
	wire v_w4719_v;
	wire v_w524_v;
	wire v_w5665_v;
	wire v_w7717_v;
	reg v_s146_v;
	wire v_w608_v;
	wire v_w6348_v;
	wire v_w7431_v;
	wire v_w2521_v;
	wire v_w383_v;
	wire v_w1958_v;
	wire v_w3584_v;
	wire v_w495_v;
	wire v_w4742_v;
	wire v_w4406_v;
	wire v_w319_v;
	wire v_w4078_v;
	wire v_w4570_v;
	wire v_w5772_v;
	wire v_w2982_v;
	wire v_w7844_v;
	wire v_w7541_v;
	wire v_w2983_v;
	wire v_w3227_v;
	wire v_w4493_v;
	wire v_w779_v;
	wire v_w25_v;
	wire v_w6116_v;
	wire v_w7069_v;
	reg v_s251_v;
	wire v_w5102_v;
	reg v_s86_v;
	wire v_w1347_v;
	wire v_w6110_v;
	reg v_s358_v;
	wire v_w5980_v;
	wire v_w4932_v;
	wire v_w3226_v;
	wire v_w7711_v;
	wire v_w6622_v;
	wire v_w6689_v;
	wire v_w8051_v;
	wire v_w3712_v;
	wire v_w519_v;
	reg v_s272_v;
	wire v_w3721_v;
	wire v_w6357_v;
	wire v_w2997_v;
	wire v_w2392_v;
	wire v_w4485_v;
	wire v_w1034_v;
	wire v_w2211_v;
	wire v_w6990_v;
	wire v_w5096_v;
	reg v_s369_v;
	wire v_w2725_v;
	wire v_w6028_v;
	wire v_w7765_v;
	wire v_w1170_v;
	wire v_w4563_v;
	wire v_w6742_v;
	wire v_w5853_v;
	wire v_w336_v;
	wire v_w4156_v;
	wire v_w2265_v;
	wire v_w1346_v;
	wire v_w7778_v;
	wire v_w4170_v;
	wire v_w373_v;
	wire v_w226_v;
	wire v_w933_v;
	wire v_w2218_v;
	wire v_w5272_v;
	wire v_w7900_v;
	wire v_w1960_v;
	wire v_w4397_v;
	wire v_w4338_v;
	wire v_w6910_v;
	reg v_s377_v;
	wire v_w7536_v;
	wire v_w7290_v;
	wire v_w2655_v;
	wire v_w3478_v;
	wire v_w1981_v;
	wire v_w1137_v;
	wire v_w720_v;
	wire v_w7889_v;
	wire v_w684_v;
	wire v_w1786_v;
	wire v_w34_v;
	wire v_w1702_v;
	wire v_w4424_v;
	wire v_w1936_v;
	wire v_w1253_v;
	wire v_w5583_v;
	wire v_w2410_v;
	wire v_w1513_v;
	wire v_w4331_v;
	reg v_s132_v;
	wire v_w2327_v;
	wire v_w5176_v;
	wire v_w3577_v;
	wire v_w7649_v;
	wire v_w4114_v;
	wire v_w3385_v;
	wire v_w4736_v;
	wire v_w6808_v;
	wire v_w5930_v;
	wire v_w7128_v;
	wire v_w1205_v;
	wire v_w5541_v;
	wire v_w3094_v;
	wire v_w549_v;
	wire v_w2924_v;
	wire v_w521_v;
	wire v_w1286_v;
	wire v_w4172_v;
	wire v_w5311_v;
	wire v_w42_v;
	wire v_w5289_v;
	reg v_s505_v;
	wire v_w7578_v;
	wire v_w3055_v;
	wire v_w6344_v;
	wire v_w7527_v;
	wire v_w3788_v;
	wire v_w4158_v;
	wire v_w7335_v;
	wire v_w4020_v;
	wire v_w3873_v;
	wire v_w1182_v;
	wire v_w5441_v;
	wire v_w8001_v;
	wire v_w1617_v;
	wire v_w6440_v;
	wire v_w8253_v;
	wire v_w4517_v;
	wire v_w11_v;
	wire v_w1996_v;
	wire v_w2690_v;
	wire v_w3239_v;
	wire v_w2661_v;
	wire v_w6183_v;
	wire v_w1852_v;
	wire v_w6355_v;
	wire v_w4703_v;
	wire v_w3291_v;
	wire v_w7708_v;
	wire v_w1569_v;
	wire v_w5751_v;
	wire v_w7209_v;
	wire v_w2090_v;
	wire v_w2662_v;
	wire v_w7032_v;
	wire v_w1697_v;
	wire v_w2772_v;
	wire v_w2992_v;
	wire v_w3481_v;
	wire v_w5083_v;
	wire v_w2756_v;
	wire v_w3701_v;
	wire v_w1540_v;
	wire v_w7721_v;
	wire v_w4909_v;
	wire v_w7739_v;
	wire v_w218_v;
	wire v_w7122_v;
	wire v_w4767_v;
	wire v_w2577_v;
	wire v_w6867_v;
	wire v_w4955_v;
	wire v_w7758_v;
	wire v_w820_v;
	wire v_w122_v;
	wire v_w6964_v;
	wire v_w3588_v;
	wire v_w5938_v;
	wire v_w2671_v;
	wire v_w4140_v;
	wire v_w3814_v;
	wire v_w1020_v;
	wire v_w7553_v;
	wire v_w3761_v;
	wire v_w7623_v;
	wire v_w6377_v;
	wire v_w3187_v;
	wire v_w932_v;
	wire v_w2239_v;
	wire v_w6757_v;
	wire v_w5911_v;
	wire v_w3463_v;
	wire v_w4979_v;
	wire v_w667_v;
	wire v_w2562_v;
	wire v_w3845_v;
	wire v_w5126_v;
	wire v_w6619_v;
	wire v_w1461_v;
	wire v_w2754_v;
	wire v_w1419_v;
	wire v_w1199_v;
	wire v_w4975_v;
	wire v_w6473_v;
	wire v_w3598_v;
	wire v_w7674_v;
	wire v_w3719_v;
	wire v_w7099_v;
	wire v_w4671_v;
	wire v_w5275_v;
	wire v_w3494_v;
	wire v_w7460_v;
	wire v_w4699_v;
	wire v_w6276_v;
	wire v_w1110_v;
	wire v_w2280_v;
	wire v_w7783_v;
	wire v_w2039_v;
	wire v_w4729_v;
	wire v_w5577_v;
	wire v_w4902_v;
	wire v_w3457_v;
	wire v_w876_v;
	wire v_w2640_v;
	wire v_w641_v;
	wire v_w2543_v;
	wire v_w5041_v;
	wire v_w1498_v;
	wire v_w3941_v;
	wire v_w7608_v;
	wire v_w6031_v;
	wire v_w6083_v;
	wire v_w7616_v;
	wire v_w6371_v;
	wire v_w7589_v;
	wire v_w7750_v;
	wire v_w1410_v;
	wire v_w6712_v;
	wire v_w2349_v;
	wire v_w7292_v;
	wire v_w3407_v;
	wire v_w6470_v;
	wire v_w3578_v;
	wire v_w1494_v;
	wire v_w3644_v;
	wire v_w4550_v;
	wire v_w5615_v;
	wire v_w7388_v;
	wire v_w4874_v;
	wire v_w5475_v;
	wire v_w4871_v;
	wire v_w7695_v;
	wire v_w2954_v;
	wire v_w2921_v;
	wire v_w5630_v;
	wire v_w4079_v;
	wire v_w1637_v;
	wire v_w7846_v;
	reg v_s168_v;
	wire v_w7594_v;
	wire v_w4184_v;
	wire v_w2182_v;
	wire v_w7584_v;
	wire v_w6252_v;
	wire v_w666_v;
	wire v_w1829_v;
	wire v_w1799_v;
	wire v_w532_v;
	wire v_w6489_v;
	wire v_w991_v;
	wire v_w1443_v;
	wire v_w6337_v;
	reg v_s40_v;
	wire v_w7443_v;
	wire v_w4027_v;
	reg v_s306_v;
	wire v_w1005_v;
	wire v_w459_v;
	wire v_w4415_v;
	wire v_w2491_v;
	reg v_s471_v;
	wire v_w7867_v;
	wire v_w5216_v;
	wire v_w986_v;
	wire v_w8240_v;
	wire v_w3957_v;
	wire v_w5810_v;
	wire v_w3952_v;
	wire v_w3058_v;
	wire v_w7848_v;
	wire v_w3639_v;
	wire v_w5483_v;
	reg v_s517_v;
	wire v_w4488_v;
	wire v_w7112_v;
	wire v_w5240_v;
	wire v_w7469_v;
	wire v_w3680_v;
	reg v_s314_v;
	wire v_w4474_v;
	wire v_w6424_v;
	wire v_w4115_v;
	wire v_w718_v;
	wire v_w5400_v;
	wire v_w4994_v;
	wire v_w3914_v;
	wire v_w7675_v;
	wire v_w5014_v;
	reg v_s244_v;
	wire v_w2752_v;
	wire v_w1147_v;
	wire v_w750_v;
	wire v_w7899_v;
	wire v_w5733_v;
	reg v_s476_v;
	wire v_w6885_v;
	wire v_w3280_v;
	wire v_w5603_v;
	wire v_w468_v;
	wire v_w2801_v;
	wire v_w456_v;
	wire v_w2988_v;
	wire v_w4181_v;
	reg v_s24_v;
	wire v_w7535_v;
	wire v_w4831_v;
	wire v_w2766_v;
	wire v_w7949_v;
	wire v_w6574_v;
	wire v_w4884_v;
	wire v_w5914_v;
	wire v_w4315_v;
	wire v_w2876_v;
	wire v_w6217_v;
	wire v_w5894_v;
	wire v_w4057_v;
	wire v_w6230_v;
	wire v_w6284_v;
	wire v_w5677_v;
	wire v_w8173_v;
	wire v_w8045_v;
	wire v_w6874_v;
	wire v_w6749_v;
	wire v_w5785_v;
	wire v_w7362_v;
	wire v_w3110_v;
	wire v_w4730_v;
	wire v_w5663_v;
	wire v_w5767_v;
	wire v_w1612_v;
	wire v_w2201_v;
	wire v_w1728_v;
	wire v_w2191_v;
	wire v_w1754_v;
	wire v_w2331_v;
	wire v_w894_v;
	wire v_w5277_v;
	wire v_w3492_v;
	wire v_w656_v;
	wire v_w4276_v;
	wire v_w4579_v;
	wire v_w2070_v;
	wire v_w702_v;
	reg v_s32_v;
	wire v_w5726_v;
	wire v_w3810_v;
	wire v_w358_v;
	wire v_w404_v;
	wire v_w4319_v;
	wire v_w6154_v;
	wire v_w3647_v;
	wire v_w4740_v;
	wire v_w1792_v;
	wire v_w939_v;
	wire v_w7718_v;
	wire v_w4271_v;
	wire v_w4988_v;
	wire v_w2872_v;
	wire v_w7053_v;
	wire v_w586_v;
	reg v_s207_v;
	wire v_w6878_v;
	wire v_w2237_v;
	wire v_w4787_v;
	wire v_w5209_v;
	wire v_w3118_v;
	wire v_w4364_v;
	wire v_w7961_v;
	wire v_w508_v;
	wire v_w6250_v;
	wire v_w1793_v;
	wire v_w6397_v;
	wire v_w6315_v;
	wire v_w7622_v;
	wire v_w1369_v;
	wire v_w4848_v;
	wire v_w3212_v;
	wire v_w6114_v;
	wire v_w4235_v;
	wire v_w1174_v;
	wire v_w1664_v;
	wire v_w4001_v;
	wire v_w578_v;
	wire v_w5291_v;
	wire v_w1662_v;
	wire v_w2590_v;
	wire v_w2346_v;
	wire v_w7954_v;
	wire v_w3306_v;
	wire v_w6049_v;
	wire v_w4088_v;
	reg v_s97_v;
	wire v_w1048_v;
	wire v_w1992_v;
	wire v_w2883_v;
	wire v_w7165_v;
	wire v_w5408_v;
	wire v_w888_v;
	wire v_w5729_v;
	wire v_w401_v;
	reg v_s309_v;
	wire v_w5178_v;
	wire v_w1812_v;
	wire v_w1003_v;
	wire v_w5290_v;
	wire v_w5039_v;
	wire v_w3354_v;
	wire v_w5943_v;
	wire v_w5018_v;
	wire v_w6155_v;
	wire v_w1072_v;
	wire v_w2172_v;
	wire v_w8061_v;
	wire v_w38_v;
	wire v_w7153_v;
	wire v_w4636_v;
	wire v_w5085_v;
	wire v_w2637_v;
	wire v_w86_v;
	wire v_w4280_v;
	wire v_w5526_v;
	wire v_w6043_v;
	wire v_w2925_v;
	wire v_w5690_v;
	wire v_w4567_v;
	wire v_w6538_v;
	wire v_w5482_v;
	wire v_w2949_v;
	wire v_w7457_v;
	wire v_w6696_v;
	reg v_s393_v;
	wire v_w3769_v;
	wire v_w4314_v;
	wire v_w3728_v;
	wire v_w4195_v;
	reg v_s479_v;
	wire v_w3008_v;
	wire v_w6581_v;
	wire v_w4546_v;
	wire v_w5399_v;
	wire v_w7477_v;
	wire v_w3591_v;
	wire v_w2019_v;
	wire v_w7656_v;
	wire v_w8226_v;
	wire v_w1983_v;
	wire v_w1736_v;
	wire v_w3742_v;
	wire v_w3004_v;
	wire v_w8136_v;
	wire v_w408_v;
	wire v_w2139_v;
	wire v_w1183_v;
	wire v_w2000_v;
	wire v_w908_v;
	wire v_w6917_v;
	wire v_w751_v;
	wire v_w52_v;
	wire v_w5699_v;
	wire v_w3670_v;
	wire v_w1471_v;
	wire v_w5215_v;
	wire v_w6394_v;
	wire v_w6836_v;
	wire v_w4138_v;
	wire v_w5877_v;
	wire v_w5586_v;
	wire v_w3822_v;
	wire v_w6903_v;
	wire v_w5817_v;
	wire v_w4588_v;
	wire v_w64_v;
	wire v_w5910_v;
	wire v_w4274_v;
	wire v_w6677_v;
	wire v_w2011_v;
	wire v_w315_v;
	wire v_w1075_v;
	wire v_w5650_v;
	wire v_w2145_v;
	wire v_w4205_v;
	reg v_s252_v;
	wire v_w1101_v;
	reg v_s461_v;
	wire v_w8066_v;
	wire v_w8129_v;
	wire v_w7706_v;
	wire v_w169_v;
	wire v_w1575_v;
	wire v_w6830_v;
	wire v_w7310_v;
	wire v_w3384_v;
	wire v_w2018_v;
	wire v_w1095_v;
	wire v_w3133_v;
	wire v_w3805_v;
	reg v_s478_v;
	wire v_w78_v;
	wire v_w6811_v;
	wire v_w6980_v;
	wire v_w6722_v;
	wire v_w4507_v;
	wire v_w7152_v;
	wire v_w2181_v;
	wire v_w452_v;
	wire v_w1912_v;
	wire v_w1660_v;
	wire v_w5682_v;
	wire v_w6816_v;
	wire v_w7777_v;
	wire v_w1337_v;
	wire v_w6495_v;
	wire v_w4377_v;
	wire v_w6324_v;
	wire v_w5725_v;
	wire v_w196_v;
	wire v_w5077_v;
	wire v_w1331_v;
	wire v_w7273_v;
	wire v_w2867_v;
	reg v_s388_v;
	reg v_s417_v;
	wire v_w1325_v;
	wire v_w4991_v;
	wire v_w7561_v;
	wire v_w569_v;
	wire v_w7086_v;
	wire v_w5940_v;
	wire v_w7028_v;
	wire v_w6531_v;
	wire v_w1502_v;
	wire v_w5515_v;
	wire v_w941_v;
	wire v_w1057_v;
	wire v_w4345_v;
	reg v_s105_v;
	reg v_s436_v;
	wire v_w4443_v;
	wire v_w6055_v;
	wire v_w372_v;
	wire v_w3727_v;
	wire v_w1824_v;
	wire v_w1354_v;
	wire v_w6267_v;
	wire v_w4270_v;
	wire v_w7127_v;
	wire v_w6071_v;
	wire v_w6795_v;
	wire v_w349_v;
	wire v_w4489_v;
	wire v_w4664_v;
	wire v_w4532_v;
	wire v_w7689_v;
	wire v_w6932_v;
	wire v_w8029_v;
	wire v_w7137_v;
	wire v_w2672_v;
	wire v_w694_v;
	reg v_s395_v;
	wire v_w7911_v;
	wire v_w5974_v;
	wire v_w8084_v;
	reg v_s13_v;
	wire v_w136_v;
	wire v_w1336_v;
	wire v_w318_v;
	wire v_w1247_v;
	wire v_w1679_v;
	wire v_w4011_v;
	wire v_w7876_v;
	wire v_w3562_v;
	wire v_w6761_v;
	wire v_w7147_v;
	wire v_o14_v;
	wire v_w4242_v;
	wire v_w8056_v;
	wire v_w6935_v;
	wire v_w1810_v;
	wire v_w3402_v;
	wire v_w1450_v;
	wire v_w2138_v;
	reg v_s6_v;
	wire v_w7145_v;
	wire v_w5652_v;
	wire v_w5826_v;
	wire v_w5567_v;
	wire v_w2121_v;
	wire v_w4135_v;
	wire v_w6341_v;
	wire v_w2023_v;
	wire v_w2670_v;
	wire v_w6320_v;
	wire v_w7898_v;
	wire v_w3642_v;
	wire v_w6229_v;
	wire v_w715_v;
	wire v_w7331_v;
	wire v_w4891_v;
	wire v_w4701_v;
	wire v_w1509_v;
	wire v_w1940_v;
	wire v_w3961_v;
	wire v_w5426_v;
	wire v_w956_v;
	wire v_w2217_v;
	wire v_w4408_v;
	wire v_w2537_v;
	wire v_w5392_v;
	wire v_w880_v;
	wire v_w1941_v;
	wire v_w2424_v;
	wire v_w341_v;
	wire v_w8206_v;
	wire v_w7253_v;
	wire v_w7078_v;
	wire v_w6978_v;
	wire v_w6467_v;
	wire v_w538_v;
	wire v_w1727_v;
	wire v_w108_v;
	wire v_w6806_v;
	wire v_w4934_v;
	wire v_w2269_v;
	wire v_w4746_v;
	wire v_w6104_v;
	wire v_w3359_v;
	wire v_w7291_v;
	wire v_w4598_v;
	wire v_w3886_v;
	wire v_w6568_v;
	wire v_w5195_v;
	wire v_w2084_v;
	wire v_w6098_v;
	reg v_s428_v;
	wire v_w5504_v;
	wire v_w7447_v;
	wire v_w3522_v;
	wire v_w7548_v;
	wire v_w7178_v;
	wire v_w7546_v;
	wire v_w6943_v;
	wire v_w6164_v;
	wire v_w2047_v;
	wire v_w1006_v;
	wire v_w2822_v;
	wire v_w5027_v;
	wire v_w4544_v;
	wire v_w5103_v;
	wire v_w2358_v;
	wire v_w1666_v;
	wire v_w6132_v;
	wire v_w3779_v;
	wire v_w1580_v;
	wire v_w7806_v;
	wire v_w6297_v;
	wire v_w7615_v;
	wire v_w2468_v;
	wire v_w4911_v;
	wire v_w8237_v;
	wire v_w7635_v;
	wire v_w7237_v;
	wire v_w3344_v;
	wire v_w3081_v;
	wire v_w1236_v;
	wire v_w1691_v;
	wire v_w5322_v;
	wire v_w7057_v;
	wire v_w6204_v;
	wire v_w2306_v;
	wire v_w727_v;
	wire v_w2510_v;
	wire v_w1078_v;
	wire v_w6308_v;
	wire v_w2683_v;
	wire v_w277_v;
	wire v_w5378_v;
	wire v_w4311_v;
	wire v_w665_v;
	wire v_w1084_v;
	reg v_s115_v;
	reg v_s5_v;
	wire v_w3128_v;
	wire v_w1856_v;
	wire v_w6376_v;
	wire v_w7268_v;
	wire v_w8134_v;
	wire v_w4505_v;
	reg v_s63_v;
	wire v_w1343_v;
	wire v_w7125_v;
	wire v_w5128_v;
	wire v_w2761_v;
	wire v_w2248_v;
	wire v_w7755_v;
	wire v_w1374_v;
	wire v_w872_v;
	wire v_w529_v;
	wire v_w307_v;
	wire v_w1466_v;
	wire v_w4606_v;
	wire v_w3357_v;
	wire v_w6019_v;
	wire v_w2817_v;
	wire v_w8044_v;
	wire v_w1599_v;
	wire v_w4087_v;
	wire v_w245_v;
	wire v_w2357_v;
	wire v_w5433_v;
	wire v_w6459_v;
	wire v_w994_v;
	wire v_w1902_v;
	wire v_w921_v;
	wire v_w7164_v;
	wire v_w3431_v;
	wire v_w2776_v;
	wire v_w613_v;
	wire v_w1281_v;
	wire v_w1000_v;
	reg v_s444_v;
	reg v_s56_v;
	wire v_w4452_v;
	wire v_w6741_v;
	wire v_w1440_v;
	wire v_w491_v;
	wire v_w2508_v;
	wire v_w1145_v;
	wire v_w1683_v;
	reg v_s405_v;
	wire v_w1307_v;
	wire v_w2732_v;
	wire v_w4250_v;
	wire v_w6680_v;
	wire v_w6636_v;
	wire v_w4450_v;
	wire v_w1726_v;
	wire v_w1254_v;
	wire v_w3029_v;
	wire v_w347_v;
	wire v_w1734_v;
	wire v_w5498_v;
	wire v_w1387_v;
	wire v_w929_v;
	wire v_w5648_v;
	wire v_w6608_v;
	wire v_w1210_v;
	wire v_w12_v;
	wire v_w2204_v;
	wire v_w3047_v;
	wire v_w7193_v;
	wire v_w1473_v;
	wire v_w8123_v;
	wire v_w7098_v;
	wire v_w2294_v;
	wire v_w3879_v;
	wire v_w7771_v;
	wire v_w935_v;
	wire v_w8002_v;
	wire v_w8097_v;
	reg v_s121_v;
	wire v_w5194_v;
	wire v_w3449_v;
	wire v_w8243_v;
	wire v_w4272_v;
	wire v_w6442_v;
	wire v_w5092_v;
	wire v_w1105_v;
	wire v_w5032_v;
	reg v_s102_v;
	wire v_w410_v;
	wire v_w4666_v;
	wire v_w8161_v;
	wire v_w6888_v;
	wire v_w2945_v;
	wire v_w6596_v;
	wire v_w1164_v;
	wire v_w7136_v;
	wire v_w7686_v;
	wire v_w6940_v;
	wire v_w4766_v;
	wire v_w4679_v;
	wire v_w5239_v;
	wire v_w4625_v;
	wire v_w2449_v;
	wire v_w1701_v;
	wire v_w1018_v;
	wire v_w3378_v;
	wire v_w522_v;
	wire v_w4704_v;
	wire v_w6454_v;
	wire v_w258_v;
	wire v_w7047_v;
	wire v_w4918_v;
	wire v_w5140_v;
	wire v_w2893_v;
	wire v_w4490_v;
	wire v_w185_v;
	wire v_w6298_v;
	wire v_w1570_v;
	wire v_w2390_v;

	assign v_w6528_v = ~(v_s355_v & v_w6499_v);
	assign v_w5688_v = ~(v_w5686_v & v_w5687_v);
	assign v_w1019_v = ~(v_w736_v & v_w1272_v);
	assign v_w4890_v = v_w3642_v ^ v_w4551_v;
	assign v_w3972_v = ~(v_w3574_v & v_w3732_v);
	assign v_w7621_v = ~(v_w1327_v & v_w7620_v);
	assign v_w7678_v = ~(v_w7078_v & v_w7677_v);
	assign v_w6429_v = v_w1424_v ^ v_w6428_v;
	assign v_w814_v = ~(v_w2300_v & v_w1299_v);
	assign v_w6766_v = ~(v_w6765_v & v_w1707_v);
	assign v_w7341_v = ~(v_w7336_v & v_w7339_v);
	assign v_w5016_v = ~(v_w2369_v & v_w2585_v);
	assign v_w3944_v = ~(v_w3732_v | v_w3943_v);
	assign v_w4594_v = ~(v_w674_v & v_s428_v);
	assign v_w5353_v = ~(v_w683_v & v_w5352_v);
	assign v_w1417_v = ~(v_w1020_v | v_w1416_v);
	assign v_w2068_v = ~(v_w8178_v);
	assign v_w7007_v = ~(v_w7006_v & v_w655_v);
	assign v_w4360_v = ~(v_w4353_v & v_w4359_v);
	assign v_w1888_v = ~(v_w1886_v & v_w1887_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s263_v<=0;
	end
	else
	begin
	v_s263_v<=v_w279_v;
	end
	end
	assign v_w3434_v = ~(v_w3095_v | v_w2620_v);
	assign v_w1243_v = ~(v_s198_v & v_w1192_v);
	assign v_w1519_v = ~(v_w1051_v & v_s234_v);
	assign v_w6954_v = ~(v_w6952_v & v_w6953_v);
	assign v_w6248_v = ~(v_w6234_v | v_w6247_v);
	assign v_w8086_v = ~(v_w6909_v | v_w6962_v);
	assign v_w1296_v = ~(v_w874_v & v_s441_v);
	assign v_w4224_v = ~(v_w4054_v & v_s330_v);
	assign v_w7289_v = ~(v_w7287_v | v_w7288_v);
	assign v_w6507_v = ~(v_w6495_v | v_w6506_v);
	assign v_w314_v = ~(v_s497_v);
	assign v_w4236_v = ~(v_w2823_v & v_s210_v);
	assign v_w7834_v = ~(v_w654_v & v_w7833_v);
	assign v_w6135_v = ~(v_w6131_v ^ v_w6134_v);
	assign v_w6143_v = ~(v_w657_v & v_s286_v);
	assign v_w5844_v = ~(v_w2137_v & v_w788_v);
	assign v_w2771_v = ~(v_w2355_v & v_s116_v);
	assign v_w3120_v = ~(v_w3108_v & v_w3119_v);
	assign v_w5487_v = ~(v_w683_v & v_w5486_v);
	assign v_w5965_v = ~(v_s270_v & v_w5786_v);
	assign v_w445_v = ~(v_w5658_v & v_w5659_v);
	assign v_w7554_v = ~(v_w7552_v & v_w7553_v);
	assign v_w1688_v = ~(v_w1419_v | v_w802_v);
	assign v_w3768_v = v_w8195_v ^ v_keyinput_92_v;
	assign v_w8160_v = ~(v_w5056_v & v_w4588_v);
	assign v_w8229_v = v_w3635_v ^ v_keyinput_113_v;
	assign v_w4354_v = ~(v_s371_v & v_w2784_v);
	assign v_w2930_v = ~(v_w2929_v);
	assign v_w5471_v = ~(v_w683_v & v_w5470_v);
	assign v_w2154_v = ~(v_w2153_v & v_w120_v);
	assign v_w121_v = ~(v_w5650_v & v_w5651_v);
	assign v_w3505_v = ~(v_w2440_v | v_w3504_v);
	assign v_w5873_v = ~(v_w5871_v & v_w5872_v);
	assign v_w7027_v = ~(v_w7025_v | v_w7026_v);
	assign v_w7211_v = ~(v_w1503_v | v_w528_v);
	assign v_w2600_v = ~(v_w2598_v | v_w2599_v);
	assign v_w6819_v = ~(v_w1412_v | v_w6571_v);
	assign v_w6346_v = ~(v_w6345_v & v_w659_v);
	assign v_w1290_v = v_s440_v ^ v_w1169_v;
	assign v_w3979_v = ~(v_w3971_v | v_w3978_v);
	assign v_w2244_v = ~(v_w2243_v);
	assign v_w7366_v = ~(v_w687_v | v_w765_v);
	assign v_w5477_v = ~(v_w5476_v | v_w4708_v);
	assign v_w6103_v = ~(v_w6077_v & v_w6080_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s19_v<=0;
	end
	else
	begin
	v_s19_v<=v_w21_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s39_v<=0;
	end
	else
	begin
	v_s39_v<=v_w46_v;
	end
	end
	assign v_w4834_v = ~(v_w2753_v | v_w2370_v);
	assign v_w3523_v = ~(v_w2827_v | v_w2833_v);
	assign v_w7525_v = ~(v_w687_v & v_w1297_v);
	assign v_w708_v = v_w2147_v & v_w2148_v;
	assign v_w5945_v = ~(v_w1624_v | v_w5734_v);
	assign v_w442_v = ~(v_w5656_v & v_w5657_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s455_v<=0;
	end
	else
	begin
	v_s455_v<=v_w508_v;
	end
	end
	assign v_w5609_v = ~(v_w5555_v & v_w5514_v);
	assign v_w4734_v = ~(v_w2342_v | v_w4733_v);
	assign v_w7244_v = ~(v_w7242_v & v_w7243_v);
	assign v_w1740_v = ~(v_w1739_v);
	assign v_w794_v = ~(v_in20_v & v_w1238_v);
	assign v_w7374_v = ~(v_w1828_v | v_w680_v);
	assign v_w6797_v = ~(v_w6788_v & v_w6796_v);
	assign v_w643_v = ~(v_w641_v | v_w642_v);
	assign v_w7229_v = ~(v_w7227_v | v_w7228_v);
	assign v_w5578_v = ~(v_s200_v & v_w676_v);
	assign v_w2127_v = ~(v_w2126_v);
	assign v_w2296_v = ~(v_w2292_v | v_w2295_v);
	assign v_w4635_v = ~(v_w674_v & v_s427_v);
	assign v_w1733_v = ~(v_w1365_v | v_w1732_v);
	assign v_w3456_v = ~(v_w3455_v ^ v_in2_v);
	assign v_w1552_v = ~(v_s271_v & v_w874_v);
	assign v_w7474_v = ~(v_w7356_v & v_w7473_v);
	assign v_w5762_v = ~(v_w5707_v & v_w1367_v);
	assign v_w1883_v = ~(v_w1384_v);
	assign v_w4446_v = ~(v_w4443_v & v_w4445_v);
	assign v_w2471_v = ~(v_w2469_v | v_w2470_v);
	assign v_w450_v = ~(v_w5765_v & v_w5768_v);
	assign v_w6544_v = ~(v_w6543_v & v_w6020_v);
	assign v_w2176_v = ~(v_w793_v & v_w2175_v);
	assign v_w6105_v = v_w1539_v ^ v_w6104_v;
	assign v_w6756_v = ~(v_w6755_v & v_w655_v);
	assign v_w612_v = v_w710_v;
	assign v_w4157_v = ~(v_w4155_v & v_w4156_v);
	assign v_w429_v = ~(v_w3371_v & v_w3378_v);
	assign v_w3415_v = ~(v_w2378_v | v_w2606_v);
	assign v_w1122_v = ~(v_w565_v & v_s38_v);
	assign v_w5283_v = ~(v_w5282_v & v_w878_v);
	assign v_w2926_v = ~(v_w2921_v | v_w2925_v);
	assign v_w1823_v = ~(v_w1632_v);
	assign v_w551_v = ~(v_w549_v | v_w550_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s488_v<=0;
	end
	else
	begin
	v_s488_v<=v_w180_v;
	end
	end
	assign v_w3073_v = ~(v_s384_v ^ v_w2655_v);
	assign v_w8222_v = v_w8221_v ^ v_keyinput_108_v;
	assign v_w3152_v = ~(v_w2607_v & v_w2833_v);
	assign v_w308_v = ~(v_w7018_v & v_w7029_v);
	assign v_w4670_v = ~(v_w4664_v & v_w4669_v);
	assign v_w5865_v = ~(v_s436_v & v_w529_v);
	assign v_w5784_v = ~(v_w2137_v & v_w602_v);
	assign v_w7556_v = ~(v_w7554_v ^ v_w7555_v);
	assign v_w2378_v = ~(v_w2374_v | v_w2377_v);
	assign v_w7097_v = ~(v_w1798_v & v_w1834_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s456_v<=0;
	end
	else
	begin
	v_s456_v<=v_w509_v;
	end
	end
	assign v_w3180_v = ~(v_w3178_v & v_w3179_v);
	assign v_w3620_v = ~(v_w3471_v & v_w3619_v);
	assign v_w7240_v = ~(v_w7237_v & v_w6578_v);
	assign v_w2259_v = ~(v_w866_v | v_w2233_v);
	assign v_w5582_v = ~(v_s119_v & v_w676_v);
	assign v_w5871_v = ~(v_w5703_v & v_w5870_v);
	assign v_w6695_v = ~(v_w6694_v & v_w6626_v);
	assign v_w628_v = ~(v_w626_v & v_w627_v);
	assign v_w4772_v = ~(v_w674_v | v_w4771_v);
	assign v_w7989_v = ~(v_s467_v | v_s363_v);
	assign v_w8178_v = v_w8177_v ^ v_keyinput_81_v;
	assign v_w8159_v = ~(v_w3992_v | v_w3993_v);
	assign v_w1371_v = ~(v_w666_v & v_s97_v);
	assign v_w2763_v = ~(v_w558_v & v_w1016_v);
	assign v_w6527_v = ~(v_w1391_v & v_w6498_v);
	assign v_w947_v = v_w946_v;
	assign v_w5932_v = ~(v_w1674_v | v_w2135_v);
	assign v_w5731_v = ~(v_w1330_v | v_w2135_v);
	assign v_w6674_v = v_w6571_v | v_w1316_v;
	assign v_w3286_v = ~(v_w2773_v | v_w2606_v);
	assign v_w224_v = ~(v_w5354_v & v_w5361_v);
	assign v_w3255_v = ~(v_w3253_v & v_w3254_v);
	assign v_w7472_v = ~(v_w7364_v & v_w7471_v);
	assign v_w5170_v = ~(v_w5168_v | v_w5169_v);
	assign v_w4709_v = ~(v_w4526_v | v_w4705_v);
	assign v_w4866_v = ~(v_w866_v & v_w4865_v);
	assign v_w6564_v = ~(v_s451_v & v_w874_v);
	assign v_w6316_v = ~(v_w6314_v & v_w6315_v);
	assign v_w2518_v = ~(v_w2516_v & v_w2517_v);
	assign v_w3722_v = ~(v_w3601_v | v_w3721_v);
	assign v_w1884_v = v_w8212_v ^ v_keyinput_103_v;
	assign v_w6147_v = ~(v_w6029_v | v_w6146_v);
	assign v_w1024_v = ~(v_in25_v | v_w1255_v);
	assign v_w6524_v = ~(v_w6522_v ^ v_w6523_v);
	assign v_w2352_v = ~(v_w991_v | v_s251_v);
	assign v_w1175_v = ~(v_s100_v | v_s398_v);
	assign v_w7662_v = ~(v_w5906_v | v_w7661_v);
	assign v_w3994_v = v_w8159_v ^ v_keyinput_66_v;
	assign v_w8028_v = ~(v_s462_v ^ v_s315_v);
	assign v_w681_v = ~(v_w2260_v | v_w2255_v);
	assign v_w1030_v = ~(v_w1032_v & v_w745_v);
	assign v_w1693_v = ~(v_w666_v & v_s101_v);
	assign v_w3197_v = ~(v_w593_v & v_s19_v);
	assign v_w1113_v = v_w8074_v ^ v_keyinput_10_v;
	assign v_w5661_v = ~(v_w420_v & v_w2738_v);
	assign v_w7266_v = ~(v_w680_v & v_w1064_v);
	assign v_w3269_v = ~(v_w2998_v ^ v_w2999_v);
	assign v_w4180_v = ~(v_w4171_v | v_w4179_v);
	assign v_w6946_v = ~(v_w6944_v | v_w6945_v);
	assign v_w7043_v = ~(v_w7036_v & v_w7042_v);
	assign v_w3715_v = ~(v_w3711_v | v_w3714_v);
	assign v_w4388_v = ~(v_w3175_v & v_w4387_v);
	assign v_w3587_v = ~(v_w2690_v);
	assign v_w463_v = ~(v_w6724_v & v_w6725_v);
	assign v_w4712_v = v_w852_v ^ v_w4414_v;
	assign v_w3922_v = v_w3801_v | v_w3918_v;
	assign v_w5842_v = ~(v_w5840_v & v_w5841_v);
	assign v_w2356_v = ~(v_w2355_v & v_s229_v);
	assign v_w1634_v = ~(v_w1616_v & v_w1633_v);
	assign v_w607_v = ~(v_w1569_v & v_w1570_v);
	assign v_w7731_v = ~(v_w1656_v | v_w1782_v);
	assign v_w425_v = ~(v_s513_v);
	assign v_w7416_v = ~(v_w679_v | v_w1834_v);
	assign v_w6120_v = ~(v_w664_v & v_s457_v);
	assign v_w3013_v = ~(v_w3012_v | v_w557_v);
	assign v_w2325_v = ~(v_w564_v & v_s248_v);
	assign v_w2819_v = ~(v_w2814_v | v_w2818_v);
	assign v_w5937_v = ~(v_w2137_v & v_w1337_v);
	assign v_w1559_v = ~(v_w1558_v & v_w613_v);
	assign v_w1315_v = ~(v_s423_v & v_w562_v);
	assign v_w5763_v = ~(v_w892_v & v_w1384_v);
	assign v_w3877_v = v_w8166_v ^ v_keyinput_71_v;
	assign v_w35_v = ~(v_w7901_v & v_w7902_v);
	assign v_w3309_v = ~(v_w2400_v | v_w2606_v);
	assign v_w2770_v = ~(v_w699_v & v_s178_v);
	assign v_w1053_v = ~(v_w1105_v & v_w1050_v);
	assign v_w6436_v = ~(v_w6434_v & v_w6435_v);
	assign v_w3435_v = ~(v_w3433_v | v_w3434_v);
	assign v_w6432_v = ~(v_w6407_v | v_w6411_v);
	assign v_w3099_v = ~(v_w3098_v & v_w2478_v);
	assign v_w5713_v = ~(v_w662_v & v_w1678_v);
	assign v_w5252_v = ~(v_w1542_v | v_w5145_v);
	assign v_w3955_v = ~(v_w3954_v & v_w3945_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s45_v<=0;
	end
	else
	begin
	v_s45_v<=v_w53_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s8_v<=0;
	end
	else
	begin
	v_s8_v<=v_w9_v;
	end
	end
	assign v_w2245_v = ~(v_w2230_v & v_w2244_v);
	assign v_w648_v = ~(v_w647_v);
	assign v_w4165_v = ~(v_w4164_v & v_w692_v);
	assign v_w1202_v = ~(v_s32_v & v_w1192_v);
	assign v_w1485_v = ~(v_w870_v & v_w1484_v);
	assign v_w6475_v = ~(v_w664_v & v_s470_v);
	assign v_w1587_v = ~(v_w1585_v | v_w1586_v);
	assign v_w4675_v = ~(v_w674_v & v_s410_v);
	assign v_w5654_v = ~(v_s107_v & v_w695_v);
	assign v_w7938_v = ~(v_w527_v & v_w1655_v);
	assign v_w3335_v = ~(v_w3333_v | v_w3334_v);
	assign v_w1165_v = ~(v_s408_v | v_w1164_v);
	assign v_w6042_v = ~(v_s477_v | v_w42_v);
	assign v_w705_v = v_w708_v & v_w709_v;
	assign v_w3832_v = ~(v_w3830_v & v_w3831_v);
	assign v_w4320_v = ~(v_w2984_v ^ v_w4319_v);
	assign v_w3028_v = ~(v_w699_v & v_s181_v);
	assign v_w6688_v = ~(v_w6684_v | v_w6687_v);
	assign v_w2338_v = ~(v_w2318_v & v_w2337_v);
	assign v_w6447_v = ~(v_w6446_v & v_w6020_v);
	assign v_w7033_v = ~(v_w1532_v | v_w6571_v);
	assign v_w5900_v = ~(v_w1602_v | v_w2135_v);
	assign v_w6362_v = ~(v_w6360_v ^ v_w6361_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s512_v<=0;
	end
	else
	begin
	v_s512_v<=v_w414_v;
	end
	end
	assign v_w2517_v = ~(v_w2484_v & v_w1131_v);
	assign v_w3017_v = ~(v_s125_v ^ v_w3016_v);
	assign v_w2659_v = v_w2658_v & v_s386_v;
	assign v_w3607_v = ~(v_w3602_v & v_w3606_v);
	assign v_w3990_v = ~(v_w3988_v & v_w3989_v);
	assign v_w7055_v = ~(v_w884_v & v_w7048_v);
	assign v_w4074_v = ~(v_w897_v & v_s262_v);
	assign v_w1919_v = ~(v_w1918_v & v_w1781_v);
	assign v_w6405_v = ~(v_w6403_v & v_w6404_v);
	assign v_w227_v = ~(v_w7717_v & v_w7718_v);
	assign v_w2519_v = v_w2515_v ^ v_w2518_v;
	assign v_w2668_v = ~(v_w2361_v | v_w2667_v);
	assign v_w1725_v = ~(v_w1723_v & v_w1724_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s273_v<=0;
	end
	else
	begin
	v_s273_v<=v_w291_v;
	end
	end
	assign v_w6372_v = ~(v_w6370_v & v_w6371_v);
	assign v_w4751_v = ~(v_w4742_v | v_w4750_v);
	assign v_w6560_v = ~(v_w6018_v | v_w1378_v);
	assign v_w1676_v = ~(v_w1673_v | v_w1675_v);
	assign v_w2617_v = ~(v_w2358_v & v_s314_v);
	assign v_w2532_v = ~(v_w2530_v & v_w2531_v);
	assign v_w3401_v = ~(v_w3023_v ^ v_w3027_v);
	assign v_w3347_v = ~(v_w3346_v & v_w1139_v);
	assign v_w4099_v = ~(v_w3160_v & v_w4098_v);
	assign v_w4854_v = ~(v_w674_v | v_w4853_v);
	assign v_w5437_v = ~(v_w5435_v | v_w5436_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s124_v<=0;
	end
	else
	begin
	v_s124_v<=v_w133_v;
	end
	end
	assign v_w5410_v = ~(v_s177_v & v_w5386_v);
	assign v_w2308_v = ~(v_w2303_v | v_w2307_v);
	assign v_w3399_v = ~(v_w3394_v | v_w3398_v);
	assign v_w5878_v = ~(v_w5876_v & v_w5877_v);
	assign v_w1082_v = ~(v_w2294_v | v_w1427_v);
	assign v_w2415_v = ~(v_w2413_v & v_w2414_v);
	assign v_w6577_v = v_w6573_v & v_w655_v;
	assign v_w1263_v = ~(v_s289_v & v_w1192_v);
	assign v_w5478_v = ~(v_w5475_v & v_w5477_v);
	assign v_w6400_v = v_s341_v ^ v_w6399_v;
	assign v_w2753_v = ~(v_w2748_v | v_w2752_v);
	assign v_w2558_v = ~(v_w2556_v & v_w2557_v);
	assign v_w4049_v = ~(v_w690_v & v_s256_v);
	assign v_w7287_v = ~(v_w687_v | v_w1734_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s449_v<=0;
	end
	else
	begin
	v_s449_v<=v_w502_v;
	end
	end
	assign v_w2345_v = v_s277_v & v_s278_v;
	assign v_w5129_v = ~(v_w5127_v | v_w5128_v);
	assign v_w5012_v = ~(v_s299_v & v_w674_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s94_v<=0;
	end
	else
	begin
	v_s94_v<=v_w102_v;
	end
	end
	assign v_w1821_v = ~(v_w1820_v & v_w1094_v);
	assign v_w454_v = ~(v_w6756_v & v_w6761_v);
	assign v_w4747_v = ~(v_w4745_v & v_w4746_v);
	assign v_w7003_v = ~(v_w1798_v & v_w1100_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s374_v<=0;
	end
	else
	begin
	v_s374_v<=v_w418_v;
	end
	end
	assign v_w6461_v = ~(v_s89_v & v_w888_v);
	assign v_w3561_v = ~(v_w1078_v | v_w3338_v);
	assign v_w2290_v = ~(v_w2289_v);
	assign v_w6733_v = ~(v_w6731_v & v_w6732_v);
	assign v_w8087_v = v_w8086_v ^ v_keyinput_17_v;
	assign v_w4065_v = ~(v_w4063_v & v_w4064_v);
	assign v_w4192_v = ~(v_w4189_v ^ v_w4191_v);
	assign v_w5628_v = ~(v_s282_v & v_w695_v);
	assign v_w7483_v = ~(v_w1418_v | v_w680_v);
	assign v_w7471_v = ~(v_w7365_v & v_w7470_v);
	assign v_w1624_v = ~(v_w1620_v | v_w1623_v);
	assign v_w3361_v = ~(v_w3126_v & v_w3360_v);
	assign v_w3353_v = ~(v_w2607_v & v_w2937_v);
	assign v_w2094_v = ~(v_w2091_v | v_w2093_v);
	assign v_w2703_v = ~(v_w2361_v | v_w2702_v);
	assign v_w4036_v = ~(v_w4035_v | v_w48_v);
	assign v_w5860_v = ~(v_w5859_v & v_w5703_v);
	assign v_w3894_v = ~(v_w3818_v & v_w3821_v);
	assign v_w1851_v = ~(v_w980_v | v_w1850_v);
	assign v_w4400_v = ~(v_w2590_v & v_w4399_v);
	assign v_w4061_v = ~(v_w185_v | v_w274_v);
	assign v_w1869_v = ~(v_w1821_v & v_w1868_v);
	assign v_w3215_v = ~(v_w3214_v & v_w3126_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s511_v<=0;
	end
	else
	begin
	v_s511_v<=v_w403_v;
	end
	end
	assign v_w7870_v = ~(v_s207_v & v_w1993_v);
	assign v_w4417_v = ~(v_w753_v | v_w4416_v);
	assign v_w2886_v = ~(v_w825_v | v_w617_v);
	assign v_w5841_v = ~(v_w662_v & v_w944_v);
	assign v_w241_v = ~(v_w5338_v & v_w5346_v);
	assign v_w2293_v = ~(v_w1192_v & v_w568_v);
	assign v_w2485_v = ~(v_w2484_v & v_w2399_v);
	assign v_w6171_v = ~(v_w6169_v & v_w6170_v);
	assign v_w3754_v = ~(v_w3735_v & v_w2706_v);
	assign v_w6011_v = ~(v_s475_v & v_w1966_v);
	assign v_w8174_v = ~(v_w4044_v | v_w4045_v);
	assign v_w5585_v = ~(v_w675_v & v_w5408_v);
	assign v_w7915_v = ~(v_s36_v & v_w6015_v);
	assign v_w8079_v = v_w6730_v & v_w6737_v;
	assign v_w48_v = ~(v_s485_v);
	assign v_w5852_v = ~(v_s343_v & v_w528_v);
	assign v_w2097_v = v_w1999_v ^ v_w1003_v;
	assign v_w3619_v = ~(v_w3617_v & v_w3618_v);
	assign v_w2339_v = ~(v_w2309_v | v_w2338_v);
	assign v_w4889_v = ~(v_w4888_v & v_w2456_v);
	assign v_w8197_v = v_w8196_v ^ v_keyinput_93_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s65_v<=0;
	end
	else
	begin
	v_s65_v<=v_w73_v;
	end
	end
	assign v_w4468_v = ~(v_w8245_v);
	assign v_w1592_v = ~(v_w1536_v & v_w1591_v);
	assign v_w6419_v = ~(v_w6418_v & v_w659_v);
	assign v_w4525_v = ~(v_w866_v | v_w556_v);
	assign v_w769_v = ~(v_w767_v | v_w768_v);
	assign v_w1595_v = ~(v_w1594_v | v_w790_v);
	assign v_w8151_v = v_w8150_v ^ v_keyinput_60_v;
	assign v_w5599_v = ~(v_w5555_v & v_w5470_v);
	assign v_w4155_v = ~(v_w2290_v & v_s294_v);
	assign v_w600_v = ~(v_w628_v & v_w2061_v);
	assign v_w6045_v = ~(v_s247_v & v_w528_v);
	assign v_w7458_v = ~(v_w1624_v & v_w680_v);
	assign v_w3723_v = ~(v_w3603_v & v_w3722_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s43_v<=0;
	end
	else
	begin
	v_s43_v<=v_w51_v;
	end
	end
	assign v_w5926_v = ~(v_w5924_v | v_w5925_v);
	assign v_w6251_v = ~(v_w6249_v & v_w6250_v);
	assign v_w1757_v = ~(v_s448_v | v_w1171_v);
	assign v_w2088_v = ~(v_w2001_v | v_w2087_v);
	assign v_w6304_v = ~(v_w6302_v & v_w6303_v);
	assign v_w5118_v = ~(v_s156_v & v_w2347_v);
	assign v_w1801_v = ~(v_w1796_v | v_w1800_v);
	assign v_w3189_v = ~(v_w2484_v & v_w3118_v);
	assign v_w322_v = ~(v_w7213_v & v_w7214_v);
	assign v_w1984_v = ~(v_w1975_v & v_w1979_v);
	assign v_w7926_v = ~(v_w527_v & v_w1026_v);
	assign v_w7701_v = ~(v_w989_v | v_w1782_v);
	assign v_w2228_v = ~(v_w2212_v | v_w2227_v);
	assign v_w2714_v = ~(v_w2478_v & v_w820_v);
	assign v_w3991_v = ~(v_w3987_v | v_w3990_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s35_v<=0;
	end
	else
	begin
	v_s35_v<=v_w41_v;
	end
	end
	assign v_w3314_v = ~(v_w3312_v & v_w3313_v);
	assign v_w397_v = ~(v_w7673_v & v_w7674_v);
	assign v_w7037_v = ~(v_w648_v ^ v_w1844_v);
	assign v_w6683_v = ~(v_w6682_v & v_w6626_v);
	assign v_w7503_v = ~(v_w7292_v | v_w7289_v);
	assign v_w5491_v = ~(v_w5489_v | v_w5490_v);
	assign v_w5619_v = ~(v_w5555_v & v_w5552_v);
	assign v_w7986_v = v_s469_v & v_s370_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s229_v<=0;
	end
	else
	begin
	v_s229_v<=v_w242_v;
	end
	end
	assign v_w4754_v = ~(v_w4753_v | v_w2342_v);
	assign v_w2041_v = v_w2039_v | v_w2040_v;
	assign v_w4330_v = v_w4326_v ^ v_w415_v;
	assign v_w7572_v = ~(v_w1870_v | v_w7571_v);
	assign v_w6569_v = ~(v_w6566_v | v_w6568_v);
	assign v_w878_v = ~(v_w876_v & v_w877_v);
	assign v_w882_v = ~(v_w686_v);
	assign v_w391_v = ~(v_w4258_v & v_w4273_v);
	assign v_w4685_v = v_w4509_v ^ v_w3632_v;
	assign v_w5825_v = ~(v_w5823_v & v_w5824_v);
	assign v_w3018_v = ~(v_w3017_v);
	assign v_w2089_v = v_w1311_v ^ v_w1997_v;
	assign v_w4644_v = ~(v_w4641_v | v_w4643_v);
	assign v_w3733_v = ~(v_w3470_v & v_w3732_v);
	assign v_w496_v = ~(v_w5702_v & v_w5711_v);
	assign v_w6791_v = ~(v_w6790_v & v_w6626_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s238_v<=0;
	end
	else
	begin
	v_s238_v<=v_w251_v;
	end
	end
	assign v_w3240_v = ~(v_w3109_v & v_w2890_v);
	assign v_w4498_v = ~(v_w3025_v | v_w1079_v);
	assign v_w6210_v = ~(v_w6187_v & v_w6190_v);
	assign v_w2144_v = ~(v_s169_v | v_s170_v);
	assign v_w4613_v = ~(v_w4611_v | v_w4612_v);
	assign v_w2492_v = ~(v_w2488_v & v_w2491_v);
	assign v_w7052_v = ~(v_w1798_v & v_w944_v);
	assign v_w5698_v = ~(v_s444_v & v_w528_v);
	assign v_w3397_v = ~(v_w2607_v & v_w2429_v);
	assign v_w2759_v = ~(v_w2754_v | v_w2758_v);
	assign v_w3293_v = ~(v_w3291_v & v_w3292_v);
	assign v_w3104_v = v_w3097_v | v_w3103_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s402_v<=0;
	end
	else
	begin
	v_s402_v<=v_w451_v;
	end
	end
	assign v_w4237_v = ~(v_w4213_v & v_w4216_v);
	assign v_w7590_v = ~(v_w7588_v & v_w7589_v);
	assign v_w4208_v = ~(v_s314_v & v_w4190_v);
	assign v_w3662_v = ~(v_w3643_v | v_w3661_v);
	assign v_w2723_v = ~(v_w558_v & v_w2722_v);
	assign v_w6130_v = ~(v_w6129_v & v_w6020_v);
	assign v_w6058_v = ~(v_w6052_v & v_w6057_v);
	assign v_w4177_v = v_w4173_v ^ v_w4176_v;
	assign v_w3468_v = ~(v_w568_v & v_w3467_v);
	assign v_w5242_v = ~(v_w5240_v | v_w5241_v);
	assign v_w928_v = ~(v_w1816_v | v_w847_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s308_v<=0;
	end
	else
	begin
	v_s308_v<=v_w331_v;
	end
	end
	assign v_w8071_v = ~(v_w554_v & v_w555_v);
	assign v_w3525_v = ~(v_w3520_v & v_w3524_v);
	assign v_w7610_v = ~(v_w1403_v & v_w1708_v);
	assign v_w4748_v = ~(v_w4589_v | v_w4741_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s29_v<=0;
	end
	else
	begin
	v_s29_v<=v_w32_v;
	end
	end
	assign v_w216_v = ~(v_w5640_v & v_w5641_v);
	assign v_w618_v = ~(v_w621_v | v_w622_v);
	assign v_w5635_v = ~(v_w420_v & v_w2585_v);
	assign v_w1542_v = ~(v_w8180_v);
	assign v_w2929_v = ~(v_s347_v ^ v_w2880_v);
	assign v_w4797_v = ~(v_w4796_v & v_w2341_v);
	assign v_w6862_v = ~(v_w1436_v | v_w1797_v);
	assign v_w332_v = ~(v_w7929_v & v_w7930_v);
	assign v_w6299_v = v_w1626_v ^ v_w6298_v;
	assign v_w1640_v = ~(v_w666_v & v_s196_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s160_v<=0;
	end
	else
	begin
	v_s160_v<=v_w169_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s78_v<=0;
	end
	else
	begin
	v_s78_v<=v_w86_v;
	end
	end
	assign v_w3362_v = ~(v_w2870_v & v_w2634_v);
	assign v_w2712_v = ~(v_w2710_v & v_w2711_v);
	assign v_w7467_v = ~(v_w7464_v | v_w7466_v);
	assign v_w961_v = ~(v_w1004_v & v_w1005_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s48_v<=0;
	end
	else
	begin
	v_s48_v<=v_w56_v;
	end
	end
	assign v_w3040_v = ~(v_w3036_v | v_w3039_v);
	assign v_w6639_v = ~(v_w6637_v & v_w6638_v);
	assign v_w7798_v = ~(v_w8128_v);
	assign v_w4173_v = v_s221_v ^ v_w4169_v;
	assign v_w6074_v = v_s271_v ^ v_w1557_v;
	assign v_w6197_v = ~(v_w6195_v & v_w6196_v);
	assign v_w5553_v = ~(v_w683_v & v_w5552_v);
	assign v_w5150_v = ~(v_w5148_v | v_w5149_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s165_v<=0;
	end
	else
	begin
	v_s165_v<=v_w174_v;
	end
	end
	assign v_w344_v = ~(v_w7201_v & v_w7202_v);
	assign v_w5790_v = ~(v_w5785_v | v_w5789_v);
	assign v_w6580_v = ~(v_w6578_v | v_w6579_v);
	assign v_w1357_v = ~(v_w666_v & v_s80_v);
	assign v_w1925_v = v_w40_v ^ v_w1924_v;
	assign v_w630_v = ~(v_w826_v);
	assign v_w3650_v = ~(v_w3649_v);
	assign v_w240_v = ~(v_w7927_v & v_w7928_v);
	assign v_w2900_v = ~(v_w565_v & v_s198_v);
	assign v_w7772_v = ~(v_w654_v & v_w7771_v);
	assign v_w1711_v = ~(v_w1373_v & v_w1384_v);
	assign v_w8111_v = ~(v_w6531_v | v_w6533_v);
	assign v_w8194_v = v_w8193_v ^ v_keyinput_91_v;
	assign v_w7505_v = ~(v_w679_v | v_w918_v);
	assign v_w3524_v = ~(v_w3522_v | v_w3523_v);
	assign v_w2936_v = ~(v_w558_v & v_w2935_v);
	assign v_w3985_v = ~(v_w3732_v & v_w2690_v);
	assign v_w7825_v = ~(v_w6642_v & v_w7660_v);
	assign v_w6458_v = v_s406_v ^ v_w6457_v;
	assign v_w1306_v = ~(v_w1304_v & v_w1305_v);
	assign v_w4136_v = ~(v_w3275_v & v_w4135_v);
	assign v_w6153_v = ~(v_w6128_v & v_w6127_v);
	assign v_w2794_v = ~(v_w2789_v | v_w2793_v);
	assign v_w428_v = ~(v_w3230_v & v_w3237_v);
	assign v_w6076_v = ~(v_w6075_v & v_w6020_v);
	assign v_w5779_v = ~(v_w5778_v & v_w5703_v);
	assign v_w1989_v = ~(v_w1975_v | v_w1988_v);
	assign v_w3109_v = ~(v_w2620_v);
	assign v_w5758_v = ~(v_w1726_v | v_w2138_v);
	assign v_w1950_v = ~(v_w1948_v & v_w1949_v);
	assign v_w7905_v = ~(v_s443_v & v_w7876_v);
	assign v_w5320_v = ~(v_w5070_v & v_w5319_v);
	assign v_w8014_v = ~(v_w8004_v & v_w8013_v);
	assign v_w5803_v = ~(v_w1355_v | v_w2135_v);
	assign v_w1755_v = ~(v_w874_v & v_s453_v);
	assign v_w5969_v = ~(v_s399_v & v_w528_v);
	assign v_w7405_v = ~(v_w8186_v);
	assign v_w3491_v = ~(v_w572_v | v_w2937_v);
	assign v_w8055_v = ~(v_w7983_v | v_w7984_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s445_v<=0;
	end
	else
	begin
	v_s445_v<=v_w498_v;
	end
	end
	assign v_w5962_v = ~(v_w662_v & v_w1834_v);
	assign v_w4930_v = ~(v_w4526_v | v_w4926_v);
	assign v_w4682_v = ~(v_w2448_v & v_w3060_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s409_v<=0;
	end
	else
	begin
	v_s409_v<=v_w458_v;
	end
	end
	assign v_w3012_v = ~(v_w3008_v | v_w3011_v);
	assign v_w6525_v = ~(v_w6524_v & v_w659_v);
	assign v_w3960_v = ~(v_w3958_v | v_w3959_v);
	assign v_w3190_v = ~(v_w558_v & v_w963_v);
	assign v_w4238_v = ~(v_w4236_v & v_w4237_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s231_v<=0;
	end
	else
	begin
	v_s231_v<=v_w244_v;
	end
	end
	assign v_w1739_v = ~(v_w918_v | v_w1337_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s144_v<=0;
	end
	else
	begin
	v_s144_v<=v_w153_v;
	end
	end
	assign v_w7614_v = ~(v_w798_v | v_w7613_v);
	assign v_w8210_v = v_w7280_v | v_w7281_v;
	assign v_w4634_v = ~(v_w4633_v & v_w673_v);
	assign v_w7671_v = v_w7669_v & v_w7670_v;
	assign v_w4698_v = ~(v_w2261_v | v_w3056_v);
	assign v_w672_v = v_w671_v;
	assign v_w6053_v = ~(v_w713_v | v_w42_v);
	assign v_w2316_v = ~(v_w565_v & v_s274_v);
	assign v_w5017_v = v_w3648_v ^ v_w4462_v;
	assign v_w1828_v = ~(v_w788_v);
	assign v_w7491_v = ~(v_w7489_v & v_w7490_v);
	assign v_w840_v = ~(v_in9_v | v_w1204_v);
	assign v_w3829_v = v_w3825_v | v_w3828_v;
	assign v_w2957_v = ~(v_w2956_v | v_w557_v);
	assign v_w7673_v = ~(v_w654_v & v_w7672_v);
	assign v_w3171_v = ~(v_w3012_v | v_w2606_v);
	assign v_w7428_v = ~(v_w7403_v & v_w7427_v);
	assign v_w5830_v = ~(v_w2137_v & v_w1401_v);
	assign v_w6082_v = ~(v_w6081_v & v_w659_v);
	assign v_w6691_v = ~(v_s414_v & v_w656_v);
	assign v_w30_v = ~(v_w7965_v & v_w7966_v);
	assign v_w5375_v = ~(v_w5371_v | v_w5374_v);
	assign v_w2962_v = ~(v_w2961_v & v_w569_v);
	assign v_w1073_v = v_w1072_v & v_w896_v;
	assign v_w4046_v = v_w8174_v ^ v_keyinput_78_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s351_v<=0;
	end
	else
	begin
	v_s351_v<=v_w389_v;
	end
	end
	assign v_w103_v = ~(v_w5660_v & v_w5661_v);
	assign v_w441_v = ~(v_w4379_v & v_w4380_v);
	assign v_w3093_v = ~(v_s28_v & v_w2355_v);
	assign v_w7169_v = ~(v_w7167_v | v_w7168_v);
	assign v_w5704_v = ~(v_w5703_v & v_w2099_v);
	assign v_w7132_v = ~(v_w528_v | v_w1925_v);
	assign v_w6063_v = ~(v_w1579_v ^ v_w6062_v);
	assign v_w2526_v = ~(v_w2308_v | v_w617_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s138_v<=0;
	end
	else
	begin
	v_s138_v<=v_w147_v;
	end
	end
	assign v_w587_v = ~(v_w827_v & v_w304_v);
	assign v_w1460_v = ~(v_w870_v & v_w1459_v);
	assign v_w8204_v = v_w5145_v | v_w1664_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s339_v<=0;
	end
	else
	begin
	v_s339_v<=v_w370_v;
	end
	end
	assign v_w1562_v = ~(v_w533_v | v_w1374_v);
	assign v_w1710_v = ~(v_w1691_v | v_w1709_v);
	assign v_w3676_v = ~(v_w3629_v | v_w3675_v);
	assign v_w5259_v = ~(v_s248_v & v_w5140_v);
	assign v_w2482_v = v_w553_v ^ v_w2481_v;
	assign v_w1896_v = ~(v_w1893_v & v_w1895_v);
	assign v_w1853_v = ~(v_w839_v);
	assign v_w1043_v = ~(v_in16_v | v_w1226_v);
	assign v_w3264_v = ~(v_s1_v | v_w404_v);
	assign v_w3043_v = ~(v_w3035_v | v_w993_v);
	assign v_w1379_v = ~(v_w1374_v | v_w1378_v);
	assign v_w8039_v = ~(v_w7991_v | v_w8038_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s122_v<=0;
	end
	else
	begin
	v_s122_v<=v_w131_v;
	end
	end
	assign v_w3632_v = ~(v_w3575_v | v_w3589_v);
	assign v_w4019_v = ~(v_w3735_v | v_w3618_v);
	assign v_w8135_v = v_w8134_v ^ v_keyinput_49_v;
	assign v_w5389_v = ~(v_w2601_v & v_w2935_v);
	assign v_w1117_v = ~(v_w809_v & v_w1354_v);
	assign v_w4279_v = ~(v_w4259_v & v_w4262_v);
	assign v_w4804_v = ~(v_w4802_v & v_w4803_v);
	assign v_w2387_v = ~(v_w2385_v & v_w2386_v);
	assign v_w305_v = ~(v_w5882_v & v_w5887_v);
	assign v_w7304_v = ~(v_w1373_v | v_w680_v);
	assign v_w5106_v = ~(v_w2461_v ^ v_w2462_v);
	assign v_w265_v = ~(v_w5150_v & v_w5151_v);
	assign v_w1759_v = ~(v_w1052_v & v_s10_v);
	assign v_w1897_v = ~(v_w1324_v | v_w1067_v);
	assign v_w6264_v = ~(v_s322_v ^ v_w6263_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s434_v<=0;
	end
	else
	begin
	v_s434_v<=v_w486_v;
	end
	end
	assign v_w5961_v = ~(v_w5703_v & v_w5960_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s83_v<=0;
	end
	else
	begin
	v_s83_v<=v_w91_v;
	end
	end
	assign v_w2541_v = ~(v_w2536_v ^ v_w2540_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s267_v<=0;
	end
	else
	begin
	v_s267_v<=v_w284_v;
	end
	end
	assign v_w8184_v = v_w8183_v ^ v_keyinput_85_v;
	assign v_w4084_v = v_w4083_v ^ v_s172_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s173_v<=0;
	end
	else
	begin
	v_s173_v<=v_w186_v;
	end
	end
	assign v_w6654_v = ~(v_s439_v & v_w656_v);
	assign v_w2530_v = ~(v_w558_v & v_w2309_v);
	assign v_w3720_v = ~(v_w3719_v | v_w1006_v);
	assign v_w1861_v = ~(v_w1642_v | v_w1656_v);
	assign v_w7773_v = ~(v_s108_v & v_w7742_v);
	assign v_w7080_v = ~(v_w7079_v & v_w655_v);
	assign v_w5429_v = ~(v_w2601_v & v_w1016_v);
	assign v_w507_v = ~(v_w6041_v & v_w6043_v);
	assign v_w7606_v = ~(v_w7605_v & v_w1438_v);
	assign v_w5870_v = ~(v_w2085_v ^ v_w2086_v);
	assign v_w6136_v = ~(v_w6135_v & v_w659_v);
	assign v_w1966_v = v_s44_v ^ v_w1965_v;
	assign v_w1333_v = ~(v_w1052_v & v_s37_v);
	assign v_w5450_v = ~(v_w5447_v & v_w5449_v);
	assign v_w175_v = ~(v_w5166_v & v_w5167_v);
	assign v_w1129_v = ~(v_w2404_v | v_w2405_v);
	assign v_w6094_v = ~(v_w6018_v | v_w1557_v);
	assign v_w60_v = v_s52_v & v_w7107_v;
	assign v_w3901_v = ~(v_w2914_v & v_w881_v);
	assign v_w7456_v = ~(v_w7442_v & v_w7445_v);
	assign v_w903_v = ~(v_w2036_v);
	assign v_w3233_v = ~(v_w3232_v & v_w3126_v);
	assign v_w6485_v = ~(v_s109_v ^ v_w6484_v);
	assign v_w475_v = ~(v_w7142_v & v_w7143_v);
	assign v_w4287_v = ~(v_w4267_v & v_w4268_v);
	assign v_w7839_v = ~(v_w1114_v & v_w7838_v);
	assign v_w4458_v = ~(v_w2803_v & v_w2618_v);
	assign v_w5356_v = ~(v_w4975_v & v_w5355_v);
	assign v_w874_v = v_w670_v;
	assign v_w4473_v = ~(v_w4471_v | v_w4472_v);
	assign v_w3648_v = ~(v_w3510_v | v_w3503_v);
	assign v_w3500_v = ~(v_w2436_v | v_w3499_v);
	assign v_w4620_v = ~(v_s434_v & v_w674_v);
	assign v_w3970_v = ~(v_w3968_v & v_w3969_v);
	assign v_w6649_v = ~(v_w1286_v | v_w1797_v);
	assign v_w7794_v = ~(v_w1783_v & v_w1119_v);
	assign v_w6018_v = ~(v_w6016_v | v_w6017_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s219_v<=0;
	end
	else
	begin
	v_s219_v<=v_w232_v;
	end
	end
	assign v_w1131_v = v_w8105_v ^ v_keyinput_29_v;
	assign v_w7306_v = ~(v_w680_v | v_w1384_v);
	assign v_w5203_v = ~(v_s90_v & v_w5141_v);
	assign v_w2878_v = ~(v_w2877_v | v_w531_v);
	assign v_w1097_v = ~(v_w2808_v | v_w2811_v);
	assign v_w7913_v = ~(v_s3_v & v_w1993_v);
	assign v_w6520_v = ~(v_w1391_v & v_w6483_v);
	assign v_w7410_v = v_w7406_v | v_w7409_v;
	assign v_w62_v = v_s54_v & v_w7107_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s400_v<=0;
	end
	else
	begin
	v_s400_v<=v_w449_v;
	end
	end
	assign v_w1526_v = ~(v_w562_v & v_s282_v);
	assign v_w3695_v = ~(v_w3513_v);
	assign v_w8069_v = v_w3126_v & v_w3315_v;
	assign v_w5883_v = ~(v_w981_v | v_w2028_v);
	assign v_w4048_v = ~(v_w692_v & v_s258_v);
	assign v_w5594_v = ~(v_s104_v & v_w676_v);
	assign v_w8148_v = v_w5878_v | v_w5881_v;
	assign v_w761_v = ~(v_w760_v);
	assign v_w8219_v = ~(v_w2387_v | v_w2390_v);
	assign v_w4971_v = ~(v_w2847_v | v_w2370_v);
	assign v_w3466_v = ~(v_w612_v & v_s4_v);
	assign v_w2187_v = ~(v_w2185_v & v_w2186_v);
	assign v_w6543_v = v_w6541_v ^ v_w6542_v;
	assign v_w2038_v = ~(v_w728_v & v_w2037_v);
	assign v_w3089_v = ~(v_w699_v & v_s188_v);
	assign v_w2112_v = ~(v_w2111_v & v_w1972_v);
	assign v_w5004_v = ~(v_w4997_v & v_w5003_v);
	assign v_w7162_v = ~(v_s396_v & v_w7113_v);
	assign v_w2263_v = ~(v_w2257_v | v_w555_v);
	assign v_w6774_v = ~(v_w1140_v & v_w1367_v);
	assign v_w3625_v = v_w3476_v ^ v_w3480_v;
	assign v_w7264_v = ~(v_w7262_v | v_w7263_v);
	assign v_w788_v = ~(v_w1132_v & v_w1133_v);
	assign v_w983_v = ~(v_w1374_v | v_w1528_v);
	assign v_w7478_v = ~(v_w7340_v & v_w7477_v);
	assign v_w2233_v = v_s170_v ^ v_w2232_v;
	assign v_w4875_v = ~(v_w2448_v & v_w2890_v);
	assign v_w4103_v = ~(v_w4102_v & v_w4093_v);
	assign v_w3129_v = ~(v_w2607_v & v_w2890_v);
	assign v_w1191_v = ~(v_s24_v & v_w562_v);
	assign v_w3674_v = ~(v_w3630_v | v_w3673_v);
	assign v_w323_v = ~(v_w7209_v & v_w7210_v);
	assign v_w7143_v = ~(v_w7118_v & v_w1313_v);
	assign v_w2285_v = ~(v_s289_v & v_w565_v);
	assign v_w6771_v = ~(v_w6770_v & v_w6626_v);
	assign v_w6588_v = ~(v_w6577_v | v_w6587_v);
	assign v_w512_v = ~(v_w6165_v & v_w6178_v);
	assign v_w3003_v = ~(v_w3001_v | v_w3002_v);
	assign v_w2594_v = v_w2587_v | v_w2593_v;
	assign v_w5197_v = ~(v_w1386_v | v_w5145_v);
	assign v_w5226_v = ~(v_w5224_v | v_w5225_v);
	assign v_w189_v = ~(v_w5403_v & v_w5409_v);
	assign v_w8120_v = ~(v_w707_v & v_w2144_v);
	assign v_w1160_v = ~(v_w1159_v & v_w377_v);
	assign v_w1997_v = ~(v_w723_v ^ v_w1065_v);
	assign v_w5580_v = ~(v_s352_v & v_w676_v);
	assign v_w5430_v = ~(v_w5428_v & v_w5429_v);
	assign v_w4247_v = ~(v_w2896_v & v_w887_v);
	assign v_w2484_v = ~(v_w993_v);
	assign v_w1647_v = ~(v_w1646_v | v_w808_v);
	assign v_w5753_v = v_w2025_v ^ v_w2026_v;
	assign v_w7804_v = ~(v_w1919_v | v_w6699_v);
	assign v_w1092_v = ~(v_w1664_v | v_w808_v);
	assign v_w1572_v = ~(v_w1051_v & v_s359_v);
	assign v_w4835_v = ~(v_w4833_v | v_w4834_v);
	assign v_w8179_v = ~(v_w1029_v ^ v_w1030_v);
	assign v_w3462_v = ~(v_in3_v & v_w3459_v);
	assign v_w5575_v = ~(v_w675_v & v_w5368_v);
	assign v_w3363_v = ~(v_w3361_v & v_w3362_v);
	assign v_w4781_v = v_w4453_v ^ v_w4496_v;
	assign v_w2809_v = ~(v_w558_v & v_w2803_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s426_v<=0;
	end
	else
	begin
	v_s426_v<=v_w477_v;
	end
	end
	assign v_w2490_v = ~(v_w2335_v | v_w538_v);
	assign v_w3409_v = ~(v_w3121_v | v_w864_v);
	assign v_w2267_v = ~(v_w793_v);
	assign v_w5318_v = ~(v_w2318_v | v_w2602_v);
	assign v_w1837_v = ~(v_w606_v);
	assign v_w4555_v = ~(v_w956_v & v_w4554_v);
	assign v_w6979_v = ~(v_w884_v & v_w6978_v);
	assign v_w2209_v = ~(v_s153_v | v_s152_v);
	assign v_w5563_v = ~(v_w675_v & v_w5320_v);
	assign v_w201_v = ~(v_w5516_v & v_w5523_v);
	assign v_w7021_v = ~(v_w1788_v & v_w944_v);
	assign v_w7544_v = ~(v_w7542_v | v_w7543_v);
	assign v_w7685_v = ~(v_w654_v & v_w7684_v);
	assign v_w7068_v = v_w1584_v ^ v_w603_v;
	assign v_w7784_v = ~(v_w654_v & v_w7783_v);
	assign v_w1013_v = ~(v_w2300_v & v_w1289_v);
	assign v_w2065_v = v_w1699_v ^ v_w894_v;
	assign v_w2194_v = ~(v_w2193_v);
	assign v_w653_v = ~(v_w1972_v & v_w7659_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s296_v<=0;
	end
	else
	begin
	v_s296_v<=v_w318_v;
	end
	end
	assign v_w6832_v = ~(v_w1020_v | v_w6579_v);
	assign v_w6282_v = ~(v_w5888_v & v_w6281_v);
	assign v_w285_v = ~(v_w7229_v & v_w7230_v);
	assign v_w2095_v = ~(v_w2092_v | v_w1297_v);
	assign v_w1909_v = ~(v_w1804_v | v_w1908_v);
	assign v_w1496_v = v_s305_v ^ v_w1150_v;
	assign v_w6384_v = ~(v_s195_v & v_w1465_v);
	assign v_w1674_v = v_s340_v ^ v_w1156_v;
	assign v_w5548_v = ~(v_s192_v & v_w5293_v);
	assign v_w5497_v = ~(v_w683_v & v_w5496_v);
	assign v_w4430_v = ~(v_w2369_v & v_w4429_v);
	assign v_w2707_v = ~(v_w558_v & v_w2706_v);
	assign v_w4575_v = ~(v_w3575_v | v_w4574_v);
	assign v_w7220_v = v_w7112_v & v_s282_v;
	assign v_w4438_v = ~(v_w4436_v | v_w4437_v);
	assign v_w5928_v = v_w631_v ^ v_w5927_v;
	assign v_w1846_v = ~(v_w1026_v);
	assign v_w6966_v = ~(v_w1101_v | v_w6608_v);
	assign v_w6775_v = ~(v_w6773_v & v_w6774_v);
	assign v_w2320_v = ~(v_w947_v | v_w531_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s217_v<=0;
	end
	else
	begin
	v_s217_v<=v_w230_v;
	end
	end
	assign v_w3567_v = ~(v_w820_v);
	assign v_w6027_v = ~(v_s158_v & v_w528_v);
	assign v_w4809_v = ~(v_w4808_v & v_w673_v);
	assign v_w6534_v = v_w8111_v ^ v_keyinput_35_v;
	assign v_w7812_v = ~(v_w1067_v | v_w1782_v);
	assign v_w4970_v = ~(v_w4968_v & v_w4969_v);
	assign v_w4367_v = ~(v_w4366_v & v_w692_v);
	assign v_w1528_v = ~(v_s283_v ^ v_w1527_v);
	assign v_w4396_v = ~(v_w4388_v | v_w4395_v);
	assign v_w4393_v = ~(v_w4392_v & v_w690_v);
	assign v_w166_v = ~(v_w5620_v & v_w5621_v);
	assign v_w6487_v = ~(v_s109_v & v_w888_v);
	assign v_w1232_v = ~(v_w1230_v & v_w1231_v);
	assign v_w1023_v = ~(v_w1249_v & v_w551_v);
	assign v_w7050_v = ~(v_w7046_v & v_w7049_v);
	assign v_w2953_v = ~(v_w2952_v & v_w697_v);
	assign v_w4130_v = ~(v_w4126_v & v_w4129_v);
	assign v_w2303_v = ~(v_w2301_v & v_w2302_v);
	assign v_w1800_v = ~(v_w1798_v & v_w1799_v);
	assign v_w3298_v = ~(v_s1_v | v_w432_v);
	assign v_w273_v = ~(v_w5556_v & v_w5557_v);
	assign v_w3137_v = ~(v_w815_v ^ v_w816_v);
	assign v_w5273_v = ~(v_w3679_v | v_w4523_v);
	assign v_w1108_v = ~(v_in11_v | v_w1210_v);
	assign v_w6486_v = ~(v_w6485_v & v_w659_v);
	assign v_w4187_v = ~(v_s221_v & v_w4169_v);
	assign v_w1394_v = ~(v_w1052_v & v_s109_v);
	assign v_w7020_v = ~(v_w6602_v | v_w7019_v);
	assign v_w6730_v = ~(v_w6729_v & v_w6626_v);
	assign v_w5571_v = ~(v_w675_v & v_w5352_v);
	assign v_w7342_v = ~(v_w680_v | v_w1866_v);
	assign v_w7029_v = ~(v_w655_v & v_w7028_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s429_v<=0;
	end
	else
	begin
	v_s429_v<=v_w480_v;
	end
	end
	assign v_w3176_v = ~(v_w3174_v & v_w3175_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s59_v<=0;
	end
	else
	begin
	v_s59_v<=v_w67_v;
	end
	end
	assign v_w5394_v = ~(v_w683_v & v_w5393_v);
	assign v_w7517_v = v_w7278_v | v_w7275_v;
	assign v_w2963_v = ~(v_w1088_v | v_w617_v);
	assign v_w730_v = ~(v_s21_v ^ v_w1179_v);
	assign v_w3791_v = ~(v_w3787_v | v_w3790_v);
	assign v_w5804_v = ~(v_w5802_v | v_w5803_v);
	assign v_w5902_v = ~(v_w892_v & v_w1837_v);
	assign v_w7843_v = ~(v_s418_v & v_w7667_v);
	assign v_w4045_v = ~(v_w690_v | v_w185_v);
	assign v_w7243_v = ~(v_w680_v & v_w1769_v);
	assign v_w4795_v = ~(v_w2343_v & v_w4794_v);
	assign v_w583_v = v_w552_v ^ v_w2964_v;
	assign v_w3404_v = ~(v_w2607_v & v_w2761_v);
	assign v_w1398_v = ~(v_w1180_v | v_w1397_v);
	assign v_w1432_v = ~(v_w1430_v & v_w1431_v);
	assign v_w1464_v = ~(v_w1463_v | v_w8_v);
	assign v_w7072_v = ~(v_w7071_v & v_w1915_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s320_v<=0;
	end
	else
	begin
	v_s320_v<=v_w346_v;
	end
	end
	assign v_w6000_v = ~(v_w662_v & v_w1453_v);
	assign v_w7088_v = v_w7081_v ^ v_w608_v;
	assign v_w5298_v = ~(v_s254_v & v_w5293_v);
	assign v_w6653_v = ~(v_w655_v & v_w6652_v);
	assign v_w1436_v = ~(v_w1435_v);
	assign v_w2092_v = ~(v_w723_v ^ v_w962_v);
	assign v_w7751_v = ~(v_w6864_v | v_w7750_v);
	assign v_w857_v = ~(v_in4_v ^ v_w1766_v);
	assign v_w2029_v = ~(v_w2014_v | v_w646_v);
	assign v_w3250_v = ~(v_w3248_v & v_w3249_v);
	assign v_w2146_v = ~(v_w2145_v);
	assign v_w7446_v = ~(v_w7442_v | v_w7445_v);
	assign v_w6944_v = ~(v_w1602_v | v_w6571_v);
	assign v_w7880_v = ~(v_w651_v & v_w7747_v);
	assign v_w3421_v = ~(v_w2568_v & v_w2566_v);
	assign v_w2162_v = ~(v_w2161_v ^ v_w176_v);
	assign v_w6650_v = v_w8187_v ^ v_keyinput_87_v;
	assign v_w3705_v = ~(v_w3493_v);
	assign v_w6266_v = ~(v_w1474_v | v_w6254_v);
	assign v_w4090_v = ~(v_w897_v & v_s255_v);
	assign v_w145_v = v_s136_v & v_w5134_v;
	assign v_w2108_v = ~(v_w2105_v | v_w2107_v);
	assign v_w2499_v = ~(v_w553_v & v_w2495_v);
	assign v_w654_v = ~(v_w652_v & v_w653_v);
	assign v_w6915_v = ~(v_w6914_v | v_w1652_v);
	assign v_w6682_v = ~(v_w6678_v ^ v_w1896_v);
	assign v_w3273_v = ~(v_w3121_v | v_w967_v);
	assign v_w6491_v = ~(v_w6457_v & v_w6463_v);
	assign v_w6921_v = ~(v_w8241_v);
	assign v_w8091_v = v_w5146_v & v_w1715_v;
	assign v_w5238_v = ~(v_w5236_v | v_w5237_v);
	assign v_w7395_v = ~(v_w7390_v & v_w7393_v);
	assign v_w8164_v = v_w8163_v ^ v_keyinput_69_v;
	assign v_w2645_v = ~(v_w2644_v | v_w387_v);
	assign v_w2789_v = v_w552_v ^ v_w2788_v;
	assign v_w110_v = ~(v_w7889_v & v_w7890_v);
	assign v_w7699_v = ~(v_s233_v & v_w7667_v);
	assign v_w3126_v = ~(v_w3125_v);
	assign v_w2540_v = v_w2539_v ^ v_w552_v;
	assign v_w1876_v = ~(v_w1874_v & v_w1875_v);
	assign v_w5561_v = ~(v_w675_v & v_w5312_v);
	assign v_w6790_v = ~(v_w1709_v ^ v_w930_v);
	assign v_w251_v = ~(v_w5322_v & v_w5328_v);
	assign v_w4691_v = ~(v_w674_v | v_w4690_v);
	assign v_w3666_v = ~(v_w3638_v | v_w3665_v);
	assign v_w5985_v = ~(v_w5693_v | v_w5984_v);
	assign v_w5365_v = ~(v_w5363_v & v_w5364_v);
	assign v_w6012_v = ~(v_w6011_v);
	assign v_w3967_v = ~(v_w3960_v & v_w3963_v);
	assign v_w4792_v = ~(v_w4781_v | v_w4528_v);
	assign v_w3288_v = ~(v_w3286_v | v_w3287_v);
	assign v_w1892_v = ~(v_w1741_v & v_w1891_v);
	assign v_w4033_v = ~(v_w2241_v | v_w2194_v);
	assign v_w5142_v = v_s8_v & v_w5141_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s347_v<=0;
	end
	else
	begin
	v_s347_v<=v_w382_v;
	end
	end
	assign v_w4381_v = ~(v_w4365_v | v_w4362_v);
	assign v_w8185_v = ~(v_w729_v | v_w680_v);
	assign v_w3160_v = ~(v_s277_v & v_w1_v);
	assign v_w5745_v = ~(v_w5740_v | v_w5744_v);
	assign v_w4633_v = ~(v_w4626_v & v_w4632_v);
	assign v_w6860_v = v_w6859_v | v_w6638_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s171_v<=0;
	end
	else
	begin
	v_s171_v<=v_w183_v;
	end
	end
	assign v_w2620_v = ~(v_w2284_v & v_w2605_v);
	assign v_w1636_v = ~(v_w875_v & v_s338_v);
	assign v_w6325_v = ~(v_w6323_v & v_w6324_v);
	assign v_w6872_v = ~(v_w6871_v);
	assign v_w7351_v = ~(v_w1125_v | v_w680_v);
	assign v_w4923_v = ~(v_w2447_v & v_w2863_v);
	assign v_w8022_v = ~(v_s460_v ^ v_s297_v);
	assign v_w2169_v = ~(v_w2168_v & v_w926_v);
	assign v_w3051_v = ~(v_w8216_v);
	assign v_w6900_v = ~(v_w1798_v & v_w1678_v);
	assign v_w3148_v = ~(v_w2639_v & v_w1124_v);
	assign v_w4240_v = ~(v_w692_v & v_w4239_v);
	assign v_w3560_v = ~(v_w3557_v & v_w3559_v);
	assign v_w160_v = v_s151_v & v_w5134_v;
	assign v_w1063_v = ~(v_w1762_v ^ v_w1769_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s497_v<=0;
	end
	else
	begin
	v_s497_v<=v_w313_v;
	end
	end
	assign v_w1032_v = ~(v_in31_v & v_w777_v);
	assign v_w2621_v = ~(v_w2619_v | v_w2620_v);
	assign v_w5001_v = ~(v_w4999_v & v_w5000_v);
	assign v_w2367_v = ~(v_w2365_v & v_w2366_v);
	assign v_w6559_v = ~(v_w5760_v & v_w6558_v);
	assign v_w2373_v = ~(v_w697_v & v_w2346_v);
	assign v_w6868_v = ~(v_w1445_v | v_w6579_v);
	assign v_w5190_v = ~(v_w5188_v | v_w5189_v);
	assign v_w4788_v = ~(v_w4786_v & v_w4787_v);
	assign v_w2384_v = v_s277_v ^ v_s278_v;
	assign v_w6418_v = ~(v_w6416_v ^ v_w6417_v);
	assign v_w6041_v = ~(v_w6036_v | v_w6040_v);
	assign v_w2579_v = ~(v_w2577_v & v_w2578_v);
	assign v_w3447_v = ~(v_s5_v & v_w2355_v);
	assign v_w214_v = ~(v_w5370_v & v_w5377_v);
	assign v_w3131_v = ~(v_w3129_v & v_w3130_v);
	assign v_w2220_v = ~(v_s131_v | v_s130_v);
	assign v_w3490_v = ~(v_w2773_v & v_w968_v);
	assign v_w3095_v = ~(v_w3091_v | v_w3094_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s322_v<=0;
	end
	else
	begin
	v_s322_v<=v_w348_v;
	end
	end
	assign v_w5915_v = ~(v_w2005_v | v_w2006_v);
	assign v_w764_v = ~(v_w762_v | v_w763_v);
	assign v_w3327_v = ~(v_w3325_v & v_w3326_v);
	assign v_w1150_v = v_w1149_v | v_s303_v;
	assign v_w7863_v = ~(v_w651_v & v_w7697_v);
	assign v_w359_v = ~(v_w4920_v & v_w4935_v);
	assign v_w3953_v = ~(v_w3566_v | v_w3735_v);
	assign v_w4124_v = ~(v_w4122_v & v_w4123_v);
	assign v_w4678_v = ~(v_w2261_v | v_w3073_v);
	assign v_w6994_v = ~(v_w6992_v | v_w6993_v);
	assign v_w3876_v = ~(v_w3872_v | v_w3875_v);
	assign v_w5401_v = ~(v_w4895_v & v_w5400_v);
	assign v_w3579_v = ~(v_w3342_v & v_w820_v);
	assign v_w2067_v = ~(v_w1373_v & v_w2066_v);
	assign v_w7079_v = ~(v_w7070_v & v_w7078_v);
	assign v_w1500_v = ~(v_w765_v & v_w1100_v);
	assign v_w4116_v = ~(v_w2306_v);
	assign v_w2276_v = ~(v_s166_v | v_s218_v);
	assign v_w6411_v = ~(v_w6409_v & v_w6410_v);
	assign v_w2200_v = ~(v_w2199_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s372_v<=0;
	end
	else
	begin
	v_s372_v<=v_w416_v;
	end
	end
	assign v_w3820_v = ~(v_w2831_v & v_w3731_v);
	assign v_w4997_v = ~(v_w4996_v & v_w866_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s101_v<=0;
	end
	else
	begin
	v_s101_v<=v_w109_v;
	end
	end
	assign v_w6822_v = ~(v_w1436_v | v_w6608_v);
	assign v_w6807_v = ~(v_w6805_v & v_w6806_v);
	assign v_w7300_v = ~(v_w7298_v | v_w7299_v);
	assign v_w2398_v = ~(v_w593_v & v_s241_v);
	assign v_w3002_v = ~(v_w2760_v ^ v_w2764_v);
	assign v_w3340_v = ~(v_s381_v & v_w693_v);
	assign v_w99_v = ~(v_w7790_v & v_w7791_v);
	assign v_w193_v = ~(v_w5434_v & v_w5443_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s155_v<=0;
	end
	else
	begin
	v_s155_v<=v_w164_v;
	end
	end
	assign v_w8212_v = v_w933_v & v_w799_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s188_v<=0;
	end
	else
	begin
	v_s188_v<=v_w201_v;
	end
	end
	assign v_w6425_v = ~(v_w6413_v | v_w6424_v);
	assign v_w1275_v = ~(v_w612_v & v_s24_v);
	assign v_w1229_v = ~(v_w1227_v & v_w1228_v);
	assign v_w780_v = ~(v_w778_v & v_w779_v);
	assign v_w4676_v = ~(v_w2265_v & v_w1124_v);
	assign v_w1169_v = v_s438_v | v_w1168_v;
	assign v_w2250_v = ~(v_s174_v | v_w2199_v);
	assign v_w5623_v = ~(v_w420_v & v_w2429_v);
	assign v_w2634_v = ~(v_w2628_v & v_w2633_v);
	assign v_w689_v = v_w4030_v | v_w885_v;
	assign v_w3103_v = v_w3102_v ^ v_w552_v;
	assign v_w1763_v = ~(v_s20_v & v_w562_v);
	assign v_w7259_v = ~(v_w680_v | v_w1003_v);
	assign v_w5589_v = ~(v_w675_v & v_w5424_v);
	assign v_w6015_v = ~(v_w527_v);
	assign v_w7470_v = ~(v_w7468_v & v_w7469_v);
	assign v_w4605_v = ~(v_w4604_v | v_w4589_v);
	assign v_w194_v = ~(v_w5444_v & v_w5451_v);
	assign v_w1945_v = ~(v_s61_v | v_s59_v);
	assign v_w1538_v = ~(v_w829_v | v_w8_v);
	assign v_w3763_v = ~(v_w3761_v & v_w3762_v);
	assign v_w2914_v = ~(v_w2910_v);
	assign v_w3753_v = ~(v_w3751_v | v_w3752_v);
	assign v_w3887_v = ~(v_w3879_v & v_w3886_v);
	assign v_w3502_v = ~(v_w3494_v & v_w3501_v);
	assign v_w2858_v = ~(v_w2848_v | v_w2857_v);
	assign v_w3918_v = ~(v_w2890_v & v_w3732_v);
	assign v_w4439_v = ~(v_w674_v & v_s429_v);
	assign v_w8060_v = ~(v_w7993_v | v_w7994_v);
	assign v_w325_v = ~(v_w7205_v & v_w7206_v);
	assign v_w7159_v = ~(v_w1378_v | v_w529_v);
	assign v_w4819_v = ~(v_w4817_v | v_w4818_v);
	assign v_w259_v = ~(v_w7856_v & v_w7857_v);
	assign v_w3875_v = ~(v_w3873_v & v_w3874_v);
	assign v_w1124_v = ~(v_w1122_v & v_w1123_v);
	assign v_w1776_v = ~(v_w8123_v);
	assign v_w2627_v = ~(v_w2246_v & v_w2626_v);
	assign v_w3496_v = v_w3495_v | v_w2238_v;
	assign v_w7340_v = v_w7336_v | v_w7339_v;
	assign v_w1761_v = ~(v_w1756_v | v_w1760_v);
	assign v_w548_v = ~(v_s219_v | v_w547_v);
	assign v_w6899_v = ~(v_w6897_v | v_w6898_v);
	assign v_w1428_v = v_s342_v ^ v_w1158_v;
	assign v_w5024_v = ~(v_w2447_v & v_w2379_v);
	assign v_w604_v = ~(v_w2162_v | v_w2192_v);
	assign v_w3232_v = v_w3051_v ^ v_w3231_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s332_v<=0;
	end
	else
	begin
	v_s332_v<=v_w360_v;
	end
	end
	assign v_w5307_v = ~(v_w5076_v | v_w5306_v);
	assign v_w4989_v = ~(v_w674_v & v_s314_v);
	assign v_w1348_v = ~(v_w1344_v | v_w1347_v);
	assign v_w6647_v = ~(v_w1749_v ^ v_w1901_v);
	assign v_w2595_v = ~(v_w580_v & v_w2594_v);
	assign v_w4245_v = ~(v_w4243_v ^ v_w4244_v);
	assign v_w2305_v = ~(v_s476_v | v_w295_v);
	assign v_w6840_v = ~(v_w1798_v & v_w1416_v);
	assign v_w1715_v = ~(v_w1053_v ^ v_w1054_v);
	assign v_w483_v = ~(v_w7138_v & v_w7139_v);
	assign v_w8108_v = ~(v_w4082_v & v_w3483_v);
	assign v_w4201_v = ~(v_w4181_v & v_w4184_v);
	assign v_w3799_v = ~(v_w3735_v | v_w2890_v);
	assign v_w4413_v = ~(v_w760_v | v_w4412_v);
	assign v_w2438_v = ~(v_w2401_v | v_w2437_v);
	assign v_w7453_v = ~(v_w7449_v | v_w7452_v);
	assign v_w7970_v = v_w8147_v ^ v_keyinput_57_v;
	assign v_w6499_v = v_w1391_v ^ v_w6498_v;
	assign v_w208_v = ~(v_w7877_v & v_w7878_v);
	assign v_w5901_v = ~(v_w5899_v | v_w5900_v);
	assign v_w4862_v = ~(v_w4860_v | v_w4861_v);
	assign v_w3800_v = ~(v_w881_v | v_w1017_v);
	assign v_w1293_v = ~(v_w1052_v & v_s443_v);
	assign v_w602_v = ~(v_w729_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s73_v<=0;
	end
	else
	begin
	v_s73_v<=v_w81_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s148_v<=0;
	end
	else
	begin
	v_s148_v<=v_w157_v;
	end
	end
	assign v_w4102_v = ~(v_w2321_v & v_s253_v);
	assign v_w6328_v = ~(v_w6029_v | v_w6327_v);
	assign v_w7668_v = ~(v_s356_v & v_w7667_v);
	assign v_w6769_v = v_w6768_v | v_w6638_v;
	assign v_w7742_v = ~(v_w654_v);
	assign v_w131_v = ~(v_w7879_v & v_w7880_v);
	assign v_w4510_v = ~(v_w3632_v | v_w4509_v);
	assign v_w7647_v = ~(v_w1190_v & v_w7646_v);
	assign v_w8167_v = v_in3_v ^ v_w3459_v;
	assign v_w7984_v = v_s470_v & v_s372_v;
	assign v_w5347_v = ~(v_s220_v & v_w5293_v);
	assign v_w5835_v = ~(v_w5834_v & v_w5703_v);
	assign v_w6162_v = ~(v_s234_v ^ v_w6161_v);
	assign v_w4907_v = ~(v_w4906_v & v_w2456_v);
	assign v_w2531_v = ~(v_w2484_v & v_w2439_v);
	assign v_w6283_v = ~(v_w6018_v | v_w1610_v);
	assign v_w7172_v = ~(v_w7117_v | v_w1405_v);
	assign v_w5847_v = ~(v_w2013_v | v_w2014_v);
	assign v_w5724_v = ~(v_w5723_v & v_w5703_v);
	assign v_w5406_v = ~(v_w4867_v | v_w5123_v);
	assign v_w3809_v = ~(v_w2847_v | v_w881_v);
	assign v_w424_v = ~(v_w3410_v & v_w3411_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s84_v<=0;
	end
	else
	begin
	v_s84_v<=v_w92_v;
	end
	end
	assign v_w1181_v = ~(v_w1172_v | v_w1180_v);
	assign v_w2295_v = ~(v_w2294_v | v_w1517_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s469_v<=0;
	end
	else
	begin
	v_s469_v<=v_w522_v;
	end
	end
	assign v_w3383_v = ~(v_w3381_v | v_w3382_v);
	assign v_w6606_v = ~(v_w6604_v | v_w6605_v);
	assign v_w4990_v = ~(v_w2265_v & v_w2803_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s301_v<=0;
	end
	else
	begin
	v_s301_v<=v_w323_v;
	end
	end
	assign v_w352_v = ~(v_w5226_v & v_w5227_v);
	assign v_w4312_v = ~(v_w2961_v | v_s364_v);
	assign v_w8075_v = v_w1246_v & v_w1247_v;
	assign v_w6392_v = ~(v_w6018_v | v_w1667_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s176_v<=0;
	end
	else
	begin
	v_s176_v<=v_w189_v;
	end
	end
	assign v_w2738_v = ~(v_w2736_v & v_w2737_v);
	assign v_w3717_v = v_w8165_v ^ v_keyinput_70_v;
	assign v_w486_v = ~(v_w4624_v & v_w4634_v);
	assign v_w6_v = ~(v_w5682_v & v_w5683_v);
	assign v_w6123_v = ~(v_w664_v & v_s458_v);
	assign v_w6751_v = ~(v_w1788_v & v_w1813_v);
	assign v_w5305_v = ~(v_s252_v & v_w5293_v);
	assign v_w4384_v = ~(v_w4383_v ^ v_s104_v);
	assign v_w4374_v = ~(v_w4372_v | v_w4373_v);
	assign v_w4056_v = v_w4054_v;
	assign v_w5655_v = ~(v_w420_v & v_w2761_v);
	assign v_w989_v = ~(v_w987_v | v_w988_v);
	assign v_w7382_v = ~(v_w7380_v | v_w7381_v);
	assign v_w6029_v = ~(v_w527_v & v_w890_v);
	assign v_w4755_v = ~(v_w4752_v | v_w4754_v);
	assign v_w5702_v = ~(v_w5700_v | v_w5701_v);
	assign v_w3601_v = ~(v_w964_v | v_w3118_v);
	assign v_w1376_v = ~(v_s398_v | v_w1375_v);
	assign v_w881_v = ~(v_w879_v & v_w880_v);
	assign v_w2973_v = ~(v_w699_v & v_s177_v);
	assign v_w7271_v = ~(v_w7269_v & v_w7270_v);
	assign v_w5557_v = ~(v_w675_v & v_w5296_v);
	assign v_w390_v = ~(v_w5580_v & v_w5581_v);
	assign v_w5168_v = ~(v_w693_v | v_w2163_v);
	assign v_w4254_v = ~(v_w4056_v & v_s332_v);
	assign v_w188_v = ~(v_w5395_v & v_w5402_v);
	assign v_w3909_v = ~(v_w3907_v | v_w3908_v);
	assign v_w879_v = ~(v_w2241_v);
	assign v_w5193_v = ~(v_w3017_v | v_w1_v);
	assign v_w111_v = ~(v_w7951_v & v_w7952_v);
	assign v_w1112_v = ~(v_w6606_v & v_w6607_v);
	assign v_w6591_v = ~(v_w1917_v & v_w655_v);
	assign v_w4110_v = ~(v_w4073_v & v_w4076_v);
	assign v_w733_v = ~(v_w710_v & v_s264_v);
	assign v_w7661_v = ~(v_w7660_v | v_w1915_v);
	assign v_w2722_v = ~(v_w2720_v & v_w2721_v);
	assign v_w6024_v = ~(v_w6014_v & v_w6023_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s345_v<=0;
	end
	else
	begin
	v_s345_v<=v_w380_v;
	end
	end
	assign v_w2287_v = ~(v_w2147_v & v_w2286_v);
	assign v_w4322_v = ~(v_w4321_v & v_w692_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s58_v<=0;
	end
	else
	begin
	v_s58_v<=v_w66_v;
	end
	end
	assign v_w8100_v = v_w5146_v & v_w1767_v;
	assign v_w6168_v = ~(v_w6166_v | v_w6167_v);
	assign v_w1278_v = ~(v_w809_v & v_w1277_v);
	assign v_w7956_v = ~(v_w527_v & v_w1725_v);
	assign v_w5108_v = ~(v_w5105_v & v_w5107_v);
	assign v_w5794_v = ~(v_w662_v & v_w1725_v);
	assign v_w7030_v = ~(v_s286_v & v_w656_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s143_v<=0;
	end
	else
	begin
	v_s143_v<=v_w152_v;
	end
	end
	assign v_w7334_v = ~(v_w679_v | v_w1445_v);
	assign v_w657_v = ~(v_w889_v);
	assign v_w7697_v = ~(v_w7024_v & v_w7696_v);
	assign v_w3903_v = ~(v_w3735_v & v_w2910_v);
	assign v_w2687_v = ~(v_w2361_v | v_w2686_v);
	assign v_w7601_v = ~(v_w1660_v | v_w7600_v);
	assign v_w4596_v = ~(v_w4594_v & v_w4595_v);
	assign v_w6703_v = ~(v_w6637_v | v_w6699_v);
	assign v_w4921_v = v_w3639_v ^ v_w4547_v;
	assign v_w6657_v = ~(v_w1065_v | v_w6579_v);
	assign v_w5948_v = ~(v_s337_v & v_w529_v);
	assign v_w6747_v = ~(v_w933_v ^ v_w799_v);
	assign v_w2834_v = ~(v_w2484_v & v_w2833_v);
	assign v_w7337_v = ~(v_w680_v | v_w1681_v);
	assign v_w5464_v = ~(v_w2369_v & v_w3060_v);
	assign v_w205_v = ~(v_w5548_v & v_w5553_v);
	assign v_w143_v = v_s134_v & v_w5134_v;
	assign v_w4095_v = ~(v_w4092_v | v_w4089_v);
	assign v_w7423_v = ~(v_w7421_v & v_w7422_v);
	assign v_w3834_v = ~(v_w2378_v & v_w3731_v);
	assign v_w4951_v = ~(v_w2447_v & v_w2833_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s386_v<=0;
	end
	else
	begin
	v_s386_v<=v_w434_v;
	end
	end
	assign v_w7655_v = ~(v_s435_v & v_w1971_v);
	assign v_w7074_v = ~(v_w7072_v & v_w7073_v);
	assign v_w5304_v = ~(v_w683_v & v_w5303_v);
	assign v_w7853_v = ~(v_w651_v & v_w7665_v);
	assign v_w5112_v = ~(v_w5100_v | v_w5111_v);
	assign v_w7820_v = ~(v_w6670_v & v_w7819_v);
	assign v_w6605_v = ~(v_w1761_v | v_w1797_v);
	assign v_w2783_v = ~(v_w531_v & v_s349_v);
	assign v_w117_v = ~(v_w7887_v & v_w7888_v);
	assign v_w2588_v = ~(v_w2585_v);
	assign v_w6616_v = ~(v_s445_v & v_w656_v);
	assign v_w2793_v = ~(v_w2790_v & v_w2792_v);
	assign v_w3668_v = ~(v_w3637_v | v_w3667_v);
	assign v_w6167_v = ~(v_w6141_v | v_w6145_v);
	assign v_w6092_v = v_w6087_v ^ v_w6091_v;
	assign v_w3557_v = ~(v_w3555_v & v_w3556_v);
	assign v_w6595_v = ~(v_w6594_v);
	assign v_w4062_v = v_w4060_v ^ v_w4061_v;
	assign v_w1355_v = v_s408_v ^ v_w1164_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s427_v<=0;
	end
	else
	begin
	v_s427_v<=v_w478_v;
	end
	end
	assign v_w1317_v = ~(v_w1316_v | v_w1180_v);
	assign v_w4912_v = ~(v_w2874_v | v_w2370_v);
	assign v_w7792_v = ~(v_w6735_v | v_w1919_v);
	assign v_w3033_v = ~(v_s104_v & v_w2355_v);
	assign v_w6575_v = ~(v_w1975_v & v_w1987_v);
	assign v_w942_v = ~(v_s368_v | v_s367_v);
	assign v_w4537_v = ~(v_w2380_v | v_w4536_v);
	assign v_w1328_v = ~(v_w1325_v & v_w1327_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s159_v<=0;
	end
	else
	begin
	v_s159_v<=v_w168_v;
	end
	end
	assign v_w6216_v = ~(v_w6184_v & v_w6183_v);
	assign v_w2565_v = v_w2564_v ^ v_w553_v;
	assign v_w2585_v = ~(v_w2583_v & v_w2584_v);
	assign v_w4182_v = ~(v_s296_v & v_w4153_v);
	assign v_w438_v = ~(v_w4809_v & v_w4816_v);
	assign v_w6478_v = ~(v_w5828_v | v_w6477_v);
	assign v_w8073_v = ~(v_w6053_v | v_w6054_v);
	assign v_w2159_v = ~(v_w2158_v | v_w531_v);
	assign v_w800_v = ~(v_w1091_v & v_w1435_v);
	assign v_w2291_v = ~(v_w2290_v & v_w569_v);
	assign v_w1879_v = ~(v_w1418_v & v_w1020_v);
	assign v_w6627_v = ~(v_w6625_v & v_w6626_v);
	assign v_w6503_v = ~(v_w5852_v & v_w6502_v);
	assign v_w912_v = ~(v_w1188_v | v_w893_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s12_v<=0;
	end
	else
	begin
	v_s12_v<=v_w13_v;
	end
	end
	assign v_w7940_v = ~(v_w527_v & v_w1126_v);
	assign v_w306_v = ~(v_w7034_v & v_w7044_v);
	assign v_w5620_v = ~(v_s157_v & v_w695_v);
	assign v_w5048_v = ~(v_w5047_v & v_w673_v);
	assign v_w7176_v = ~(v_w7117_v | v_w1427_v);
	assign v_w778_v = v_w1174_v & v_w1175_v;
	assign v_w815_v = ~(v_w3068_v ^ v_w3080_v);
	assign v_w2658_v = v_w2657_v & v_s385_v;
	assign v_w5996_v = ~(v_w5994_v & v_w5995_v);
	assign v_w7451_v = ~(v_w687_v | v_w1135_v);
	assign v_w1579_v = v_w1578_v ^ v_s265_v;
	assign v_w7452_v = ~(v_w7450_v | v_w7451_v);
	assign v_w1811_v = ~(v_w1351_v & v_w1734_v);
	assign v_w5629_v = ~(v_w420_v & v_w2439_v);
	assign v_w1969_v = ~(v_w1968_v);
	assign v_w5549_v = ~(v_w3468_v | v_w2602_v);
	assign v_w506_v = ~(v_w1147_v & v_w6596_v);
	assign v_w3534_v = ~(v_w3530_v & v_w3533_v);
	assign v_w3645_v = ~(v_w3523_v | v_w3526_v);
	assign v_w10_v = ~(v_w7911_v & v_w7912_v);
	assign v_w5405_v = ~(v_w4865_v | v_w5404_v);
	assign v_w3781_v = ~(v_w2773_v | v_w881_v);
	assign v_w8036_v = ~(v_w7994_v | v_w8035_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s16_v<=0;
	end
	else
	begin
	v_s16_v<=v_w17_v;
	end
	end
	assign v_w417_v = ~(v_w5652_v & v_w5653_v);
	assign v_w7481_v = ~(v_w7479_v & v_w7480_v);
	assign v_w4277_v = ~(v_w2883_v ^ v_s362_v);
	assign v_w6734_v = ~(v_w1727_v | v_w797_v);
	assign v_w4144_v = ~(v_w4136_v | v_w4143_v);
	assign v_w6848_v = ~(v_w656_v | v_w6847_v);
	assign v_w7004_v = ~(v_w7002_v & v_w7003_v);
	assign v_w3863_v = ~(v_w3735_v | v_w2399_v);
	assign v_w5720_v = ~(v_w5718_v & v_w5719_v);
	assign v_w1557_v = ~(v_s268_v ^ v_w1556_v);
	assign v_w8015_v = ~(v_w8003_v & v_w8014_v);
	assign v_w140_v = v_s131_v & v_w5134_v;
	assign v_w2647_v = ~(v_w2646_v | v_w401_v);
	assign v_w3083_v = ~(v_w2484_v & v_w3077_v);
	assign v_w2855_v = ~(v_w2294_v | v_w1628_v);
	assign v_w7272_v = v_w7268_v | v_w7271_v;
	assign v_w5211_v = ~(v_s161_v & v_w5140_v);
	assign v_w1218_v = ~(v_s99_v & v_w1192_v);
	assign v_w5035_v = ~(v_w5034_v | v_w2457_v);
	assign v_w5849_v = ~(v_w5693_v | v_w5848_v);
	assign v_w3839_v = ~(v_w3837_v & v_w3838_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s74_v<=0;
	end
	else
	begin
	v_s74_v<=v_w82_v;
	end
	end
	assign v_w1924_v = ~(v_w999_v | v_w8_v);
	assign v_w3529_v = ~(v_w3526_v | v_w3528_v);
	assign v_w3760_v = v_w3756_v | v_w3759_v;
	assign v_w7732_v = ~(v_w6927_v | v_w7731_v);
	assign v_w6871_v = v_w1663_v ^ v_w6870_v;
	assign v_w6794_v = ~(v_w6792_v | v_w6793_v);
	assign v_w1437_v = ~(v_w1091_v);
	assign v_w4043_v = ~(v_w4041_v & v_w4042_v);
	assign v_w6897_v = ~(v_w6602_v | v_w6896_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s452_v<=0;
	end
	else
	begin
	v_s452_v<=v_w505_v;
	end
	end
	assign v_w1140_v = ~(v_w6571_v);
	assign v_w1459_v = ~(v_s339_v ^ v_w1155_v);
	assign v_w596_v = ~(v_w594_v | v_w595_v);
	assign v_w4942_v = ~(v_w4941_v | v_w4528_v);
	assign v_w671_v = ~(v_w889_v & v_w890_v);
	assign v_w4524_v = v_w3679_v ^ v_w4523_v;
	assign v_w1807_v = ~(v_w1286_v | v_w1806_v);
	assign v_w3238_v = ~(v_s1_v | v_w387_v);
	assign v_w5555_v = ~(v_w2245_v | v_w5554_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s460_v<=0;
	end
	else
	begin
	v_s460_v<=v_w513_v;
	end
	end
	assign v_w2781_v = ~(v_w2780_v & v_s349_v);
	assign v_w5505_v = ~(v_w5503_v | v_w5504_v);
	assign v_w770_v = ~(v_w1108_v | v_w1057_v);
	assign v_w4617_v = ~(v_w4616_v | v_w2264_v);
	assign v_w4198_v = ~(v_w4196_v | v_w4197_v);
	assign v_w4947_v = ~(v_w3647_v | v_w4545_v);
	assign v_w6145_v = ~(v_w1528_v ^ v_w6144_v);
	assign v_w4368_v = ~(v_w8243_v);
	assign v_w7983_v = ~(v_s470_v | v_s372_v);
	assign v_w4785_v = ~(v_w4784_v & v_w673_v);
	assign v_w4936_v = v_s329_v & v_w674_v;
	assign v_w5869_v = ~(v_w5867_v | v_w5868_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s37_v<=0;
	end
	else
	begin
	v_s37_v<=v_w44_v;
	end
	end
	assign v_w1062_v = v_w710_v & v_in33_v;
	assign v_w260_v = ~(v_w5790_v & v_w5792_v);
	assign v_w5019_v = ~(v_w878_v & v_w4538_v);
	assign v_w968_v = ~(v_w967_v);
	assign v_w7352_v = ~(v_w7350_v | v_w7351_v);
	assign v_w1382_v = ~(v_w1379_v | v_w1381_v);
	assign v_w7842_v = v_w8081_v ^ v_keyinput_14_v;
	assign v_w1188_v = ~(v_w1187_v);
	assign v_w4434_v = ~(v_w4433_v & v_w2343_v);
	assign v_w219_v = ~(v_w7723_v & v_w7724_v);
	assign v_w8031_v = ~(v_s463_v ^ v_s317_v);
	assign v_w832_v = ~(v_w1515_v & v_w1516_v);
	assign v_w430_v = ~(v_w3147_v & v_w3148_v);
	assign v_w2272_v = ~(v_w2271_v & v_s250_v);
	assign v_w6620_v = ~(v_w6595_v & v_w6619_v);
	assign v_w1865_v = ~(v_w1863_v & v_w1864_v);
	assign v_w4653_v = ~(v_w4646_v & v_w4652_v);
	assign v_w1549_v = ~(v_w665_v & v_s245_v);
	assign v_w2718_v = ~(v_s382_v ^ v_w2653_v);
	assign v_w2279_v = ~(v_w2277_v & v_w2278_v);
	assign v_w4387_v = ~(v_s395_v & v_w4054_v);
	assign v_w2697_v = ~(v_w2693_v | v_w2696_v);
	assign v_w712_v = ~(v_w711_v | v_s312_v);
	assign v_w5658_v = ~(v_s396_v & v_w695_v);
	assign v_w5742_v = ~(v_w5741_v & v_w5703_v);
	assign v_w5554_v = ~(v_w2597_v & v_w681_v);
	assign v_w3906_v = ~(v_w3902_v | v_w3905_v);
	assign v_w7433_v = ~(v_w7386_v & v_w7432_v);
	assign v_w3929_v = ~(v_w3927_v & v_w3928_v);
	assign v_w5562_v = ~(v_s241_v & v_w676_v);
	assign v_w5467_v = ~(v_w5465_v | v_w5466_v);
	assign v_w4825_v = v_w968_v ^ v_w4408_v;
	assign v_w2418_v = ~(v_w2416_v | v_w2417_v);
	assign v_w8156_v = ~(v_w1078_v | v_w2602_v);
	assign v_w1116_v = ~(v_s43_v & v_w562_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s131_v<=0;
	end
	else
	begin
	v_s131_v<=v_w140_v;
	end
	end
	assign v_w6511_v = ~(v_w1391_v & v_w6489_v);
	assign v_w7645_v = v_w1966_v & v_w7644_v;
	assign v_w385_v = ~(v_w5202_v & v_w5203_v);
	assign v_w3582_v = ~(v_w3060_v | v_w852_v);
	assign v_w4337_v = ~(v_s116_v ^ v_w4326_v);
	assign v_w8027_v = ~(v_w7999_v | v_w8026_v);
	assign v_w5319_v = ~(v_w5317_v | v_w5318_v);
	assign v_w4539_v = ~(v_w3509_v & v_w4538_v);
	assign v_w5744_v = ~(v_w5742_v & v_w5743_v);
	assign v_w1192_v = ~(v_w710_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s421_v<=0;
	end
	else
	begin
	v_s421_v<=v_w472_v;
	end
	end
	assign v_w7329_v = ~(v_w7327_v | v_w7328_v);
	assign v_w6737_v = ~(v_w6733_v | v_w6736_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s233_v<=0;
	end
	else
	begin
	v_s233_v<=v_w246_v;
	end
	end
	assign v_w7579_v = ~(v_w1709_v | v_w7578_v);
	assign v_w6379_v = v_w1667_v ^ v_w6378_v;
	assign v_w509_v = ~(v_w6084_v & v_w6095_v);
	assign v_w5568_v = ~(v_s229_v & v_w676_v);
	assign v_w2473_v = ~(v_w2439_v | v_w2309_v);
	assign v_w6281_v = ~(v_w664_v & v_s463_v);
	assign v_w1767_v = ~(v_w856_v ^ v_w857_v);
	assign v_w1605_v = ~(v_w874_v & v_s322_v);
	assign v_w5110_v = ~(v_w4525_v & v_w5106_v);
	assign v_w1228_v = ~(v_w612_v & v_s373_v);
	assign v_w4574_v = ~(v_w4572_v | v_w4573_v);
	assign v_w6801_v = ~(v_w6799_v | v_w6800_v);
	assign v_w1773_v = v_s7_v & v_w960_v;
	assign v_w6623_v = ~(v_w6618_v | v_w6622_v);
	assign v_w5645_v = ~(v_w420_v & v_w2937_v);
	assign v_w5529_v = ~(v_w5527_v & v_w5528_v);
	assign v_w5547_v = ~(v_w683_v & v_w5546_v);
	assign v_w1009_v = ~(v_w2755_v & v_w2757_v);
	assign v_w3034_v = ~(v_w3032_v & v_w3033_v);
	assign v_w6950_v = ~(v_w6592_v & v_w1853_v);
	assign v_w723_v = ~(v_w722_v);
	assign v_w6208_v = ~(v_w5686_v & v_w6207_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s170_v<=0;
	end
	else
	begin
	v_s170_v<=v_w182_v;
	end
	end
	assign v_w5422_v = ~(v_w5420_v & v_w5421_v);
	assign v_w754_v = ~(v_w753_v);
	assign v_w6587_v = ~(v_w6586_v | v_w6579_v);
	assign v_w4843_v = v_w4457_v ^ v_w4555_v;
	assign v_w7869_v = ~(v_w651_v & v_w7716_v);
	assign v_w5771_v = ~(v_w5769_v | v_w5770_v);
	assign v_w6484_v = v_w1391_v ^ v_w6483_v;
	assign v_w6684_v = ~(v_w6681_v & v_w6683_v);
	assign v_w8038_v = ~(v_w7992_v | v_w8037_v);
	assign v_w5992_v = ~(v_w5990_v | v_w5991_v);
	assign v_w3305_v = ~(v_w3109_v & v_w2690_v);
	assign v_w7495_v = ~(v_w7317_v & v_w7494_v);
	assign v_w6829_v = v_w6824_v ^ v_w802_v;
	assign v_w4999_v = ~(v_w4998_v & v_w878_v);
	assign v_w278_v = ~(v_w5115_v & v_w5116_v);
	assign v_w4558_v = ~(v_w4456_v & v_w4557_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s162_v<=0;
	end
	else
	begin
	v_s162_v<=v_w171_v;
	end
	end
	assign v_w7435_v = ~(v_w7371_v | v_w7368_v);
	assign v_w1626_v = ~(v_s320_v ^ v_w1625_v);
	assign v_w5264_v = ~(v_s172_v & v_s1_v);
	assign v_w3249_v = ~(v_w2922_v & v_w2634_v);
	assign v_w6686_v = ~(v_w1798_v & v_w1309_v);
	assign v_w790_v = v_w788_v ^ v_w789_v;
	assign v_w2001_v = ~(v_w2000_v | v_w1323_v);
	assign v_w7234_v = ~(v_s264_v & v_w7113_v);
	assign v_w3732_v = ~(v_w3731_v);
	assign v_w395_v = ~(v_w7852_v & v_w7853_v);
	assign v_w759_v = ~(v_w757_v & v_w758_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s416_v<=0;
	end
	else
	begin
	v_s416_v<=v_w467_v;
	end
	end
	assign v_w2592_v = ~(v_w2589_v | v_w2591_v);
	assign v_w1677_v = ~(v_w1052_v & v_s122_v);
	assign v_w5084_v = ~(v_w8192_v);
	assign v_w1864_v = ~(v_w1125_v & v_w1096_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s52_v<=0;
	end
	else
	begin
	v_s52_v<=v_w60_v;
	end
	end
	assign v_w4363_v = ~(v_w2756_v | v_s106_v);
	assign v_w1615_v = ~(v_w1606_v & v_w839_v);
	assign v_w2307_v = ~(v_w2306_v | v_w568_v);
	assign v_w4067_v = ~(v_w2330_v ^ v_s262_v);
	assign v_w2198_v = ~(v_w2195_v & v_w2197_v);
	assign v_w7714_v = ~(v_w6968_v | v_w7713_v);
	assign v_w701_v = v_w700_v | v_w531_v;
	assign v_w2360_v = ~(v_w2356_v & v_w2359_v);
	assign v_w4150_v = ~(v_w690_v & v_w4149_v);
	assign v_w1252_v = ~(v_w1250_v & v_w1251_v);
	assign v_w59_v = v_s51_v & v_w7107_v;
	assign v_w5261_v = ~(v_w5145_v | v_w1582_v);
	assign v_w7816_v = ~(v_s416_v & v_w7667_v);
	assign v_w2417_v = ~(v_w2331_v);
	assign v_w2773_v = ~(v_w2769_v | v_w2772_v);
	assign v_w866_v = v_w865_v;
	assign v_w698_v = ~(v_w2354_v | v_w544_v);
	assign v_w6020_v = ~(v_w1786_v | v_w658_v);
	assign v_w3631_v = ~(v_w3582_v | v_w3588_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s33_v<=0;
	end
	else
	begin
	v_s33_v<=v_w37_v;
	end
	end
	assign v_w2230_v = ~(v_w2200_v & v_w2229_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s46_v<=0;
	end
	else
	begin
	v_s46_v<=v_w54_v;
	end
	end
	assign v_w3405_v = ~(v_w3109_v & v_w3338_v);
	assign v_w4467_v = ~(v_w2575_v | v_w2585_v);
	assign v_w2529_v = v_w2528_v ^ v_w552_v;
	assign v_w7160_v = ~(v_w7117_v | v_w1380_v);
	assign v_w7293_v = ~(v_w7289_v & v_w7292_v);
	assign v_w5281_v = ~(v_w3612_v | v_w5280_v);
	assign v_w4141_v = ~(v_w4140_v & v_w692_v);
	assign v_w3765_v = ~(v_w3142_v & v_w881_v);
	assign v_w2033_v = v_w1135_v | v_w2032_v;
	assign v_w8142_v = ~(v_w6637_v | v_w6768_v);
	assign v_w4053_v = ~(v_w4039_v | v_w4052_v);
	assign v_w150_v = v_s141_v & v_w5134_v;
	assign v_w3217_v = ~(v_w2607_v & v_w3216_v);
	assign v_w6563_v = ~(v_w6552_v | v_w6562_v);
	assign v_w7199_v = ~(v_w1610_v | v_w528_v);
	assign v_w6758_v = ~(v_w6592_v & v_w997_v);
	assign v_w7022_v = ~(v_w1798_v & v_w788_v);
	assign v_w4461_v = ~(v_w2379_v | v_w2297_v);
	assign v_w7849_v = ~(v_w6570_v & v_w7848_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s473_v<=0;
	end
	else
	begin
	v_s473_v<=v_w526_v;
	end
	end
	assign v_w1933_v = ~(v_w1926_v & v_w1932_v);
	assign v_w2583_v = ~(v_w2579_v | v_w2582_v);
	assign v_w1870_v = ~(v_w1454_v & v_w1682_v);
	assign v_w16_v = ~(v_w5616_v & v_w5617_v);
	assign v_w6446_v = ~(v_s354_v ^ v_w6445_v);
	assign v_w5700_v = ~(v_w5698_v & v_w5699_v);
	assign v_w2525_v = ~(v_w2487_v | v_w2524_v);
	assign v_w2678_v = ~(v_w558_v & v_w2671_v);
	assign v_w7422_v = ~(v_w608_v & v_w680_v);
	assign v_w3030_v = ~(v_w3028_v & v_w3029_v);
	assign v_w7036_v = ~(v_w6639_v & v_w7035_v);
	assign v_w2429_v = ~(v_w2416_v);
	assign v_w6743_v = ~(v_w6592_v & v_w1119_v);
	assign v_w4321_v = v_s117_v ^ v_w4320_v;
	assign v_w900_v = ~(v_w1681_v ^ v_w1999_v);
	assign v_w6967_v = ~(v_w6965_v | v_w6966_v);
	assign v_w1154_v = v_w1153_v | v_s323_v;
	assign v_w7562_v = ~(v_w1653_v & v_w7561_v);
	assign v_w738_v = ~(v_w740_v | v_w741_v);
	assign v_w2251_v = v_w2249_v | v_w2250_v;
	assign v_w6196_v = ~(v_w657_v & v_s304_v);
	assign v_w7170_v = ~(v_s107_v & v_w7113_v);
	assign v_w386_v = ~(v_w3242_v & v_w3252_v);
	assign v_w1312_v = ~(v_w1311_v | v_w1064_v);
	assign v_w680_v = ~(v_w679_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s361_v<=0;
	end
	else
	begin
	v_s361_v<=v_w402_v;
	end
	end
	assign v_w674_v = ~(v_w673_v);
	assign v_w5210_v = ~(v_w5208_v | v_w5209_v);
	assign v_w5090_v = ~(v_w674_v & v_s266_v);
	assign v_w6884_v = ~(v_w6882_v | v_w6883_v);
	assign v_w1858_v = ~(v_w1855_v & v_w1857_v);
	assign v_w1611_v = v_w1374_v | v_w1610_v;
	assign v_w1937_v = ~(v_s64_v | v_s63_v);
	assign v_w1203_v = ~(v_w612_v & v_s423_v);
	assign v_w4480_v = ~(v_w3641_v | v_w4479_v);
	assign v_w5445_v = ~(v_w4863_v | v_w4773_v);
	assign v_w316_v = v_w2299_v | v_w2477_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s319_v<=0;
	end
	else
	begin
	v_s319_v<=v_w344_v;
	end
	end
	assign v_w6481_v = ~(v_s89_v & v_w6457_v);
	assign v_w7131_v = ~(v_s29_v & v_w7113_v);
	assign v_w4651_v = ~(v_w4642_v | v_w4589_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s376_v<=0;
	end
	else
	begin
	v_s376_v<=v_w420_v;
	end
	end
	assign v_w4642_v = v_w1008_v ^ v_w4514_v;
	assign v_w2976_v = v_s361_v ^ v_w2647_v;
	assign v_w7006_v = ~(v_w6997_v & v_w7005_v);
	assign v_w1282_v = ~(v_w1279_v & v_w1281_v);
	assign v_w619_v = v_w3062_v ^ v_w553_v;
	assign v_w3870_v = ~(v_w3862_v & v_w3869_v);
	assign v_w4487_v = ~(v_w2967_v | v_w2965_v);
	assign v_w1712_v = ~(v_w1707_v & v_w1711_v);
	assign v_w4879_v = ~(v_w4878_v & v_w673_v);
	assign v_w236_v = ~(v_w7711_v & v_w7712_v);
	assign v_w2511_v = ~(v_w2509_v | v_w2510_v);
	assign v_w289_v = ~(v_w7067_v & v_w7080_v);
	assign v_w1208_v = ~(v_s76_v & v_w1192_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s178_v<=0;
	end
	else
	begin
	v_s178_v<=v_w191_v;
	end
	end
	assign v_w6841_v = ~(v_w6839_v & v_w6840_v);
	assign v_w4995_v = v_w4399_v ^ v_w2575_v;
	assign v_w5581_v = ~(v_w675_v & v_w5393_v);
	assign v_w7325_v = v_w7321_v | v_w7324_v;
	assign v_w1489_v = ~(v_w588_v | v_w8_v);
	assign v_w4531_v = v_w963_v ^ v_w4420_v;
	assign v_w6072_v = ~(v_s86_v & v_w6055_v);
	assign v_w6368_v = ~(v_w6363_v & v_w6367_v);
	assign v_w637_v = ~(v_w2940_v);
	assign v_w6809_v = ~(v_w6808_v & v_w6626_v);
	assign v_w2445_v = v_w2383_v ^ v_w2444_v;
	assign v_w7194_v = ~(v_s333_v & v_w7112_v);
	assign v_w3602_v = ~(v_w3598_v & v_w1006_v);
	assign v_w945_v = ~(v_w944_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s317_v<=0;
	end
	else
	begin
	v_s317_v<=v_w342_v;
	end
	end
	assign v_w5638_v = ~(v_s318_v & v_w695_v);
	assign v_w2343_v = ~(v_w2342_v);
	assign v_w2694_v = ~(v_w558_v & v_w755_v);
	assign v_w822_v = ~(v_w2300_v & v_w1715_v);
	assign v_w3444_v = ~(v_w2976_v & v_w2634_v);
	assign v_w4269_v = v_w4267_v ^ v_w4268_v;
	assign v_w6908_v = ~(v_w6906_v & v_w6907_v);
	assign v_w7828_v = ~(v_s442_v & v_w7667_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s300_v<=0;
	end
	else
	begin
	v_s300_v<=v_w322_v;
	end
	end
	assign v_w1525_v = ~(v_w809_v & v_w1524_v);
	assign v_w3442_v = ~(v_w3440_v & v_w3441_v);
	assign v_w3551_v = ~(v_w3490_v & v_w3550_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s119_v<=0;
	end
	else
	begin
	v_s119_v<=v_w128_v;
	end
	end
	assign v_w6991_v = ~(v_w6592_v & v_w766_v);
	assign v_w4225_v = ~(v_w4223_v & v_w4224_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s75_v<=0;
	end
	else
	begin
	v_s75_v<=v_w83_v;
	end
	end
	assign v_w2241_v = v_w2240_v ^ v_w181_v;
	assign v_w6546_v = ~(v_w657_v | v_w6545_v);
	assign v_w6393_v = ~(v_w6391_v | v_w6392_v);
	assign v_w4905_v = ~(v_w4902_v | v_w4904_v);
	assign v_w7274_v = ~(v_w1324_v & v_w680_v);
	assign v_w5164_v = ~(v_w693_v | v_w2162_v);
	assign v_w3312_v = ~(v_s278_v & v_w693_v);
	assign v_w4013_v = ~(v_w4012_v & v_w3732_v);
	assign v_w1418_v = ~(v_w1416_v);
	assign v_w4650_v = ~(v_w4648_v & v_w4649_v);
	assign v_w5100_v = ~(v_w5096_v & v_w5099_v);
	assign v_w7232_v = ~(v_w7117_v | v_w1582_v);
	assign v_w6704_v = ~(v_w6702_v | v_w6703_v);
	assign v_w3818_v = ~(v_w3816_v & v_w3817_v);
	assign v_w7333_v = v_w7329_v | v_w7332_v;
	assign v_w7248_v = ~(v_w7246_v & v_w7247_v);
	assign v_w6593_v = ~(v_w6592_v & v_w1769_v);
	assign v_w8078_v = v_w8077_v ^ v_keyinput_12_v;
	assign v_w8218_v = v_w8217_v ^ v_keyinput_106_v;
	assign v_w2441_v = ~(v_w2392_v | v_w2440_v);
	assign v_w2638_v = ~(v_w2263_v & v_w2600_v);
	assign v_w3628_v = ~(v_w3573_v);
	assign v_w5689_v = ~(v_w662_v & v_w788_v);
	assign v_w5293_v = ~(v_w683_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s298_v<=0;
	end
	else
	begin
	v_s298_v<=v_w320_v;
	end
	end
	assign v_w6526_v = ~(v_s400_v ^ v_w1700_v);
	assign v_w1344_v = ~(v_w1343_v | v_w1180_v);
	assign v_w1245_v = ~(v_w1243_v & v_w1244_v);
	assign v_w6726_v = ~(v_w656_v & v_s409_v);
	assign v_w4959_v = ~(v_w4957_v | v_w4958_v);
	assign v_w6492_v = ~(v_w6464_v & v_w6466_v);
	assign v_w3945_v = ~(v_w1078_v & v_w3732_v);
	assign v_w4656_v = ~(v_w3629_v ^ v_w4575_v);
	assign v_w760_v = ~(v_w821_v & v_w822_v);
	assign v_w6125_v = ~(v_w1539_v & v_w6098_v);
	assign v_w4697_v = ~(v_w4695_v & v_w4696_v);
	assign v_w286_v = ~(v_w7225_v & v_w7226_v);
	assign v_w3605_v = ~(v_w3603_v & v_w3604_v);
	assign v_w7851_v = ~(v_w7742_v & v_s420_v);
	assign v_o18_v = v_w8010_v ^ v_w8011_v;
	assign v_w7494_v = ~(v_w7318_v & v_w7493_v);
	assign v_w5071_v = ~(v_w5062_v & v_w5070_v);
	assign v_w2171_v = ~(v_w2170_v & v_w181_v);
	assign v_w1744_v = ~(v_w1338_v & v_w1743_v);
	assign v_w4313_v = ~(v_w4293_v | v_w4294_v);
	assign v_w3248_v = ~(v_w3126_v & v_w3247_v);
	assign v_w7787_v = ~(v_w998_v | v_w1782_v);
	assign v_w4154_v = v_s296_v ^ v_w4153_v;
	assign v_w2102_v = ~(v_w1910_v | v_w1804_v);
	assign v_w4283_v = ~(v_w4276_v & v_w4282_v);
	assign v_w4304_v = ~(v_w4300_v & v_w4303_v);
	assign v_w7929_v = ~(v_s309_v & v_w6015_v);
	assign v_w5971_v = ~(v_w5707_v & v_w1696_v);
	assign v_w6570_v = v_w6569_v | v_w1800_v;
	assign v_w3074_v = ~(v_w2361_v | v_w3073_v);
	assign v_w435_v = ~(v_w2673_v & v_w3123_v);
	assign v_w2546_v = ~(v_w2536_v | v_w2540_v);
	assign v_w1171_v = ~(v_w497_v & v_w1170_v);
	assign v_w7631_v = ~(v_w7630_v & v_w7240_v);
	assign v_w2216_v = ~(v_s141_v | v_s143_v);
	assign v_w7744_v = ~(v_w6871_v | v_w1919_v);
	assign v_w1397_v = v_s343_v ^ v_w1160_v;
	assign v_w4750_v = ~(v_w4743_v & v_w4749_v);
	assign v_w4472_v = ~(v_w2833_v | v_w2831_v);
	assign v_w6157_v = ~(v_w6156_v & v_w6020_v);
	assign v_w3804_v = ~(v_w3802_v | v_w3803_v);
	assign v_w2504_v = v_w2503_v ^ v_w552_v;
	assign v_w3563_v = ~(v_w3561_v | v_w3562_v);
	assign v_w7357_v = ~(v_w7352_v & v_w7355_v);
	assign v_w2165_v = v_w295_v & v_w2150_v;
	assign v_w1274_v = ~(v_s14_v & v_w1192_v);
	assign v_w5808_v = ~(v_s339_v & v_w529_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s373_v<=0;
	end
	else
	begin
	v_s373_v<=v_w417_v;
	end
	end
	assign v_w7123_v = ~(v_w7118_v & v_w1767_v);
	assign v_w4089_v = v_s253_v ^ v_w2321_v;
	assign v_w4230_v = ~(v_w4226_v | v_w4229_v);
	assign v_w3419_v = ~(v_w2635_v | v_w2363_v);
	assign v_w4042_v = ~(v_w692_v & v_w274_v);
	assign v_w4762_v = ~(v_w4761_v & v_w878_v);
	assign v_w632_v = ~(v_w634_v & v_w635_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s401_v<=0;
	end
	else
	begin
	v_s401_v<=v_w450_v;
	end
	end
	assign v_w5141_v = ~(v_w8153_v);
	assign v_w135_v = v_s126_v & v_w5134_v;
	assign v_w3158_v = ~(v_w3156_v | v_w3157_v);
	assign v_w5105_v = ~(v_w5104_v & v_w878_v);
	assign v_w5381_v = ~(v_w5379_v | v_w5380_v);
	assign v_w1132_v = ~(v_w1508_v | v_w1511_v);
	assign v_w1859_v = ~(v_w1650_v | v_w1655_v);
	assign v_w7882_v = ~(v_w651_v & v_w7753_v);
	assign v_w5768_v = ~(v_w5767_v & v_w2113_v);
	assign v_w7814_v = ~(v_w6688_v & v_w7813_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s480_v<=0;
	end
	else
	begin
	v_s480_v<=v_w18_v;
	end
	end
	assign v_w6655_v = v_w6571_v | v_w1302_v;
	assign v_w5600_v = ~(v_s77_v & v_w676_v);
	assign v_w6428_v = ~(v_w6426_v & v_w6427_v);
	assign v_w1241_v = ~(v_w612_v & v_s193_v);
	assign v_w18_v = ~(v_w7116_v & v_w7119_v);
	assign v_w5811_v = v_w5810_v ^ v_w632_v;
	assign v_w1223_v = ~(v_w1221_v & v_w1222_v);
	assign v_w6700_v = ~(v_w6638_v | v_w6699_v);
	assign v_w6488_v = ~(v_w657_v & v_s355_v);
	assign v_w2505_v = ~(v_w2500_v ^ v_w2504_v);
	assign v_w3741_v = v_w3737_v | v_w3740_v;
	assign v_w7258_v = ~(v_w7249_v & v_w7257_v);
	assign v_w4227_v = ~(v_w2823_v & v_s316_v);
	assign v_w239_v = ~(v_w7864_v & v_w7865_v);
	assign v_w2887_v = ~(v_w2875_v | v_w2886_v);
	assign v_w5286_v = ~(v_w8155_v);
	assign v_w243_v = ~(v_w5329_v & v_w5337_v);
	assign v_w995_v = ~(v_w1018_v & v_w1019_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s234_v<=0;
	end
	else
	begin
	v_s234_v<=v_w247_v;
	end
	end
	assign v_w661_v = ~(v_w2122_v & v_w2105_v);
	assign v_w3063_v = ~(v_w618_v | v_w619_v);
	assign v_w3568_v = ~(v_w3567_v & v_w2722_v);
	assign v_w890_v = ~(v_w1190_v);
	assign v_w8057_v = ~(v_w7987_v | v_w7988_v);
	assign v_w5348_v = ~(v_w5007_v & v_w5126_v);
	assign v_w6226_v = v_w1490_v ^ v_w6225_v;
	assign v_w4106_v = ~(v_w4100_v & v_w4105_v);
	assign v_w6271_v = ~(v_w6269_v & v_w6270_v);
	assign v_w6919_v = ~(v_w6592_v & v_w1650_v);
	assign v_w1139_v = ~(v_w1137_v | v_w1138_v);
	assign v_w1238_v = ~(v_w1236_v & v_w1237_v);
	assign v_w387_v = ~(v_s508_v);
	assign v_w7810_v = ~(v_w6679_v);
	assign v_w5393_v = ~(v_w4913_v & v_w5392_v);
	assign v_w3743_v = ~(v_w3732_v | v_w3118_v);
	assign v_w8063_v = v_w866_v ^ v_w4391_v;
	assign v_w473_v = ~(v_w5488_v & v_w5497_v);
	assign v_w576_v = ~(v_w1546_v | v_w1547_v);
	assign v_w6084_v = ~(v_w6070_v | v_w6083_v);
	assign v_w6455_v = ~(v_s354_v & v_w6445_v);
	assign v_w757_v = ~(v_w858_v ^ v_w859_v);
	assign v_w7067_v = ~(v_w7065_v | v_w7066_v);
	assign v_w3736_v = ~(v_w3735_v | v_w3485_v);
	assign v_w2232_v = ~(v_w531_v | v_w707_v);
	assign v_w5649_v = ~(v_w420_v & v_w2967_v);
	assign v_w420_v = ~(v_w695_v);
	assign v_w1556_v = ~(v_w1555_v | v_w8_v);
	assign v_w5591_v = ~(v_w675_v & v_w5432_v);
	assign v_w2231_v = ~(v_w955_v | v_w531_v);
	assign v_w109_v = ~(v_w7778_v & v_w7779_v);
	assign v_w2829_v = ~(v_w2820_v | v_w2828_v);
	assign v_w978_v = ~(v_w976_v | v_w977_v);
	assign v_w304_v = ~(v_s496_v);
	assign v_w5934_v = v_w1351_v ^ v_w2078_v;
	assign v_w5532_v = ~(v_w4591_v & v_w5531_v);
	assign v_w2106_v = ~(v_w1914_v | v_w1996_v);
	assign v_w591_v = ~(v_w589_v | v_w590_v);
	assign v_w818_v = ~(v_w565_v & v_s82_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s135_v<=0;
	end
	else
	begin
	v_s135_v<=v_w144_v;
	end
	end
	assign v_w4064_v = ~(v_w887_v & v_w897_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s41_v<=0;
	end
	else
	begin
	v_s41_v<=v_w49_v;
	end
	end
	assign v_w5598_v = ~(v_s83_v & v_w676_v);
	assign v_w1237_v = ~(v_w612_v & v_s120_v);
	assign v_w1294_v = ~(v_w1292_v & v_w1293_v);
	assign v_w2166_v = v_w185_v & v_w2144_v;
	assign v_w4267_v = ~(v_w4265_v | v_w4266_v);
	assign v_w813_v = ~(v_w565_v & v_s27_v);
	assign v_w5397_v = ~(v_w2601_v & v_w1017_v);
	assign v_w5427_v = ~(v_w4805_v | v_w5123_v);
	assign v_w2557_v = ~(v_w565_v & v_s227_v);
	assign v_w5385_v = ~(v_w683_v & v_w5384_v);
	assign v_w6381_v = ~(v_w6350_v | v_w6380_v);
	assign v_w1804_v = ~(v_w1188_v | v_w1803_v);
	assign v_w739_v = ~(v_w737_v | v_w738_v);
	assign v_w2882_v = ~(v_w2881_v | v_w531_v);
	assign v_w4133_v = ~(v_w4131_v | v_w4132_v);
	assign v_w4405_v = ~(v_w2935_v | v_w4404_v);
	assign v_w4169_v = ~(v_w2571_v);
	assign v_w4291_v = ~(v_w2884_v & v_s362_v);
	assign v_w3704_v = ~(v_w3692_v | v_w3703_v);
	assign v_w481_v = ~(v_w5270_v & v_w5288_v);
	assign v_w4584_v = ~(v_w4583_v ^ v_w3679_v);
	assign v_w3626_v = ~(v_w3603_v & v_w3595_v);
	assign v_w5991_v = ~(v_w1286_v | v_w2138_v);
	assign v_w7307_v = ~(v_w679_v | v_w1813_v);
	assign v_w4647_v = ~(v_w8252_v);
	assign v_w4764_v = ~(v_w2369_v & v_w2738_v);
	assign v_w53_v = v_s45_v & v_w7107_v;
	assign v_w4877_v = ~(v_w4868_v | v_w4876_v);
	assign v_w7871_v = ~(v_w651_v & v_w7722_v);
	assign v_w7317_v = v_w7313_v | v_w7316_v;
	assign v_w7745_v = ~(v_w1094_v | v_w1782_v);
	assign v_w7884_v = ~(v_w651_v & v_w7759_v);
	assign v_w5718_v = ~(v_w5703_v & v_w5717_v);
	assign v_w4552_v = ~(v_w4551_v | v_w3643_v);
	assign v_w3984_v = ~(v_w3760_v & v_w3983_v);
	assign v_w130_v = ~(v_w7748_v & v_w7749_v);
	assign v_w1654_v = ~(v_w1634_v & v_w1653_v);
	assign v_w1349_v = ~(v_w666_v & v_s75_v);
	assign v_w455_v = ~(v_w6820_v & v_w6833_v);
	assign v_w7663_v = ~(v_w606_v | v_w1782_v);
	assign v_w1943_v = ~(v_w1941_v & v_w1942_v);
	assign v_w6996_v = ~(v_w6995_v);
	assign v_w1652_v = ~(v_w1624_v | v_w1632_v);
	assign v_w170_v = ~(v_w7943_v & v_w7944_v);
	assign v_w5236_v = ~(v_w1488_v | v_w5145_v);
	assign v_w6589_v = ~(v_s452_v & v_w656_v);
	assign v_w8244_v = v_w4466_v | v_w4467_v;
	assign v_w1054_v = ~(v_in13_v ^ v_w1217_v);
	assign v_w835_v = ~(v_w1488_v | v_w808_v);
	assign v_w5756_v = ~(v_w5754_v | v_w5755_v);
	assign v_w4433_v = v_w3480_v ^ v_w4422_v;
	assign v_w7941_v = ~(v_s123_v & v_w2143_v);
	assign v_w7746_v = ~(v_w7744_v | v_w7745_v);
	assign v_w777_v = ~(v_w775_v & v_w776_v);
	assign v_w153_v = v_s144_v & v_w5134_v;
	assign v_w3292_v = ~(v_w2749_v & v_w2634_v);
	assign v_w5905_v = v_w607_v & v_w606_v;
	assign v_w4556_v = ~(v_w4457_v & v_w4555_v);
	assign v_w3853_v = ~(v_w3845_v & v_w3852_v);
	assign v_w3070_v = ~(v_w699_v & v_s185_v);
	assign v_w6586_v = ~(v_w6585_v);
	assign v_w3888_v = ~(v_w3878_v | v_w3887_v);
	assign v_w1195_v = ~(v_w1193_v & v_w1194_v);
	assign v_w4176_v = ~(v_w4174_v & v_w4175_v);
	assign v_w4449_v = ~(v_w851_v & v_w3060_v);
	assign v_w4037_v = ~(v_w4029_v | v_w4036_v);
	assign v_w1760_v = ~(v_w1758_v & v_w1759_v);
	assign v_w7684_v = ~(v_w7054_v & v_w7683_v);
	assign v_w1010_v = ~(v_w1386_v | v_w2294_v);
	assign v_w296_v = ~(v_w3166_v & v_w3170_v);
	assign v_w4661_v = ~(v_w4589_v | v_w4660_v);
	assign v_w2432_v = v_w2418_v | v_w2431_v;
	assign v_w8182_v = v_w3369_v & v_w881_v;
	assign v_w6752_v = ~(v_w1798_v & v_w1362_v);
	assign v_w3932_v = ~(v_w3558_v | v_w3735_v);
	assign v_w5959_v = ~(v_w5957_v & v_w5958_v);
	assign v_w5545_v = ~(v_w5037_v & v_w4433_v);
	assign v_w3380_v = ~(v_w2607_v & v_w2863_v);
	assign v_w5075_v = ~(v_w2265_v & v_w2317_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s260_v<=0;
	end
	else
	begin
	v_s260_v<=v_w276_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s430_v<=0;
	end
	else
	begin
	v_s430_v<=v_w481_v;
	end
	end
	assign v_w6881_v = ~(v_w884_v & v_w6872_v);
	assign v_w1077_v = ~(v_w2294_v | v_w1380_v);
	assign v_w4465_v = ~(v_w4463_v | v_w4464_v);
	assign v_w5109_v = ~(v_w5103_v | v_w5108_v);
	assign v_w4162_v = ~(v_w4137_v & v_w4139_v);
	assign v_w5714_v = ~(v_w2137_v & v_w1435_v);
	assign v_w2375_v = ~(v_w2355_v & v_s231_v);
	assign v_w4323_v = ~(v_w4317_v & v_w4322_v);
	assign v_w915_v = v_w1080_v & v_w908_v;
	assign v_w2806_v = ~(v_w2804_v & v_w2805_v);
	assign v_w1918_v = v_w883_v ^ v_keyinput_6_v;
	assign v_w5136_v = ~(v_s163_v | v_w5135_v);
	assign v_w1176_v = ~(v_s44_v | v_s79_v);
	assign v_w1134_v = ~(v_w1482_v | v_w1486_v);
	assign v_w6865_v = ~(v_w6637_v | v_w6859_v);
	assign v_w1794_v = ~(v_w666_v & v_s419_v);
	assign v_w3613_v = ~(v_w3610_v | v_w3612_v);
	assign v_w7753_v = ~(v_w7751_v & v_w7752_v);
	assign v_w725_v = ~(v_w1825_v | v_w1858_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s329_v<=0;
	end
	else
	begin
	v_s329_v<=v_w357_v;
	end
	end
	assign v_w1868_v = ~(v_w1865_v & v_w1867_v);
	assign v_w2013_v = ~(v_w2012_v | v_w1026_v);
	assign v_w4431_v = ~(v_w3452_v | v_w4430_v);
	assign v_w2630_v = ~(v_w2455_v & v_w2248_v);
	assign v_w1766_v = ~(v_w1764_v & v_w1765_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s134_v<=0;
	end
	else
	begin
	v_s134_v<=v_w143_v;
	end
	end
	assign v_w1287_v = ~(v_w1286_v);
	assign v_w5368_v = ~(v_w4972_v & v_w5367_v);
	assign v_w1915_v = ~(v_w1913_v & v_w1914_v);
	assign v_w500_v = ~(v_w7907_v & v_w7908_v);
	assign v_w6335_v = ~(v_w664_v & v_s465_v);
	assign v_w5080_v = ~(v_w5076_v | v_w5079_v);
	assign v_w6641_v = ~(v_w656_v | v_w6640_v);
	assign v_w1213_v = ~(v_w1211_v & v_w1212_v);
	assign v_w4735_v = ~(v_w4732_v | v_w4734_v);
	assign v_w5778_v = ~(v_w5776_v ^ v_w5777_v);
	assign v_w2597_v = ~(v_w2247_v | v_w2251_v);
	assign v_w1873_v = ~(v_w800_v & v_w1438_v);
	assign v_w298_v = ~(v_w5074_v & v_w5075_v);
	assign v_w1703_v = ~(v_w1044_v ^ v_w1273_v);
	assign v_w834_v = ~(v_w832_v | v_w833_v);
	assign v_w7260_v = ~(v_w687_v | v_w1287_v);
	assign v_w552_v = ~(v_w2454_v & v_w556_v);
	assign v_w3565_v = ~(v_w3338_v & v_w1078_v);
	assign v_w4021_v = ~(v_w3733_v & v_w4020_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s350_v<=0;
	end
	else
	begin
	v_s350_v<=v_w388_v;
	end
	end
	assign v_w327_v = ~(v_w7007_v & v_w7012_v);
	assign v_w2852_v = ~(v_w2851_v);
	assign v_w6456_v = ~(v_w6454_v & v_w6455_v);
	assign v_w662_v = ~(v_w660_v | v_w661_v);
	assign v_w4356_v = ~(v_w4354_v & v_w4355_v);
	assign v_w4071_v = ~(v_s261_v & v_w693_v);
	assign v_w6750_v = ~(v_w6748_v & v_w6749_v);
	assign v_w2093_v = v_w1902_v ^ v_w2092_v;
	assign v_w1511_v = ~(v_w1509_v & v_w1510_v);
	assign v_w4545_v = ~(v_w3523_v | v_w4544_v);
	assign v_w7449_v = ~(v_w7447_v | v_w7448_v);
	assign v_w8195_v = v_w3735_v & v_w2738_v;
	assign v_w23_v = ~(v_w7122_v & v_w7123_v);
	assign v_w6242_v = ~(v_w1490_v & v_w6211_v);
	assign v_w639_v = v_w2839_v | v_w2859_v;
	assign v_w3307_v = ~(v_w3301_v | v_w3306_v);
	assign v_w819_v = ~(v_w2300_v & v_w1354_v);
	assign v_w141_v = v_s132_v & v_w5134_v;
	assign v_w2470_v = ~(v_w2399_v | v_w2317_v);
	assign v_w1120_v = ~(v_s14_v & v_w564_v);
	assign v_w2321_v = v_s249_v ^ v_w2320_v;
	assign v_w1501_v = ~(v_s298_v & v_w562_v);
	assign v_w5499_v = ~(v_w872_v | v_w2370_v);
	assign v_w2843_v = ~(v_w2841_v & v_w2842_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s202_v<=0;
	end
	else
	begin
	v_s202_v<=v_w215_v;
	end
	end
	assign v_w4305_v = ~(v_w692_v & v_w4304_v);
	assign v_w3381_v = ~(v_w3379_v & v_w3380_v);
	assign v_w4813_v = ~(v_w2347_v & v_w2749_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s50_v<=0;
	end
	else
	begin
	v_s50_v<=v_w58_v;
	end
	end
	assign v_w1304_v = ~(v_w874_v & v_s439_v);
	assign v_w7011_v = ~(v_w1507_v | v_w6571_v);
	assign v_w1184_v = ~(v_w1182_v & v_w1183_v);
	assign v_w1297_v = ~(v_w1295_v & v_w1296_v);
	assign v_w3049_v = v_w2741_v & v_w2744_v;
	assign v_w1187_v = ~(v_w1185_v & v_w1186_v);
	assign v_w5796_v = ~(v_w1351_v | v_w2138_v);
	assign v_w464_v = ~(v_w7897_v & v_w7898_v);
	assign v_w7501_v = ~(v_w7499_v | v_w7500_v);
	assign v_w469_v = ~(v_w7842_v & v_w7843_v);
	assign v_w3538_v = ~(v_w3536_v | v_w3537_v);
	assign v_w8093_v = v_w6141_v ^ v_w6145_v;
	assign v_w3493_v = ~(v_w3491_v | v_w3492_v);
	assign v_w5608_v = ~(v_s33_v & v_w676_v);
	assign v_w1224_v = ~(v_s110_v & v_w1192_v);
	assign v_w1512_v = ~(v_w989_v | v_w788_v);
	assign v_w7829_v = ~(v_w6619_v);
	assign v_w1488_v = ~(v_w1259_v ^ v_w739_v);
	assign v_w847_v = ~(v_w845_v | v_w846_v);
	assign v_w3756_v = ~(v_w3754_v & v_w3755_v);
	assign v_w1625_v = v_w721_v & v_s7_v;
	assign v_w7972_v = ~(v_w527_v & v_w1187_v);
	assign v_w2076_v = ~(v_w1342_v ^ v_w722_v);
	assign v_w6744_v = ~(v_w1714_v ^ v_w799_v);
	assign v_w7767_v = ~(v_s88_v & v_w7742_v);
	assign v_w6768_v = ~(v_w6766_v ^ v_w6767_v);
	assign v_w4566_v = ~(v_w3561_v | v_w4565_v);
	assign v_w1455_v = ~(v_w1052_v & v_s195_v);
	assign v_w1507_v = v_s303_v ^ v_w1149_v;
	assign v_w3263_v = ~(v_w3261_v | v_w3262_v);
	assign v_w4823_v = ~(v_w4822_v | v_w4528_v);
	assign v_w2126_v = ~(v_w1782_v | v_w1918_v);
	assign v_w3997_v = v_w873_v & v_w881_v;
	assign v_w4731_v = ~(v_w4729_v | v_w4730_v);
	assign v_w5188_v = ~(v_w1380_v | v_w5145_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s181_v<=0;
	end
	else
	begin
	v_s181_v<=v_w194_v;
	end
	end
	assign v_w6934_v = ~(v_w6931_v & v_w6933_v);
	assign v_w3933_v = ~(v_w3931_v | v_w3932_v);
	assign v_w4627_v = v_w4447_v ^ v_w4580_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s316_v<=0;
	end
	else
	begin
	v_s316_v<=v_w341_v;
	end
	end
	assign v_w946_v = ~(v_s173_v | v_s172_v);
	assign v_w282_v = ~(v_w7233_v & v_w7234_v);
	assign v_w7537_v = ~(v_w7535_v & v_w7536_v);
	assign v_w2667_v = ~(v_s386_v ^ v_w2658_v);
	assign v_w926_v = ~(v_w924_v & v_w925_v);
	assign v_w4869_v = v_w958_v ^ v_w4553_v;
	assign v_w635_v = v_w2052_v | v_w1642_v;
	assign v_w3151_v = ~(v_s1_v | v_w355_v);
	assign v_w7332_v = v_w7330_v | v_w7331_v;
	assign v_w3609_v = ~(v_w3600_v & v_w3608_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s338_v<=0;
	end
	else
	begin
	v_s338_v<=v_w369_v;
	end
	end
	assign v_w934_v = v_w1287_v ^ v_w1003_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s501_v<=0;
	end
	else
	begin
	v_s501_v<=v_w354_v;
	end
	end
	assign v_w3793_v = ~(v_w3731_v & v_w1088_v);
	assign v_w6678_v = ~(v_w1328_v);
	assign v_w2791_v = ~(v_w2773_v);
	assign v_w6032_v = ~(v_w6030_v | v_w6031_v);
	assign v_w1029_v = v_in30_v ^ v_w1271_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s220_v<=0;
	end
	else
	begin
	v_s220_v<=v_w233_v;
	end
	end
	assign v_w7064_v = ~(v_w1140_v & v_s270_v);
	assign v_w735_v = ~(v_w796_v | v_w969_v);
	assign v_w3367_v = ~(v_s383_v & v_w693_v);
	assign v_w4324_v = ~(v_w4311_v | v_w4323_v);
	assign v_w6864_v = ~(v_w6855_v & v_w6863_v);
	assign v_w8190_v = v_w8189_v ^ v_keyinput_89_v;
	assign v_w3455_v = ~(v_w3453_v & v_w3454_v);
	assign v_w4564_v = ~(v_w4452_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s201_v<=0;
	end
	else
	begin
	v_s201_v<=v_w214_v;
	end
	end
	assign v_w3691_v = ~(v_w3543_v);
	assign v_w5309_v = ~(v_w5307_v & v_w5308_v);
	assign v_w2333_v = ~(v_w569_v | v_w2332_v);
	assign v_w3780_v = ~(v_w3778_v | v_w3779_v);
	assign v_w5734_v = ~(v_w662_v);
	assign v_w2131_v = ~(v_w2108_v);
	assign v_w7864_v = ~(v_s226_v & v_w1993_v);
	assign v_w2578_v = ~(v_w2358_v & v_s299_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s315_v<=0;
	end
	else
	begin
	v_s315_v<=v_w340_v;
	end
	end
	assign v_w534_v = ~(v_w1577_v & v_w1581_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s243_v<=0;
	end
	else
	begin
	v_s243_v<=v_w256_v;
	end
	end
	assign v_w4931_v = ~(v_w4929_v | v_w4930_v);
	assign v_w27_v = ~(v_w7126_v & v_w7127_v);
	assign v_w419_v = ~(v_w7169_v & v_w7170_v);
	assign v_w7936_v = ~(v_w527_v & v_w1824_v);
	assign v_w2709_v = v_w553_v ^ v_w2708_v;
	assign v_w6982_v = ~(v_w6980_v & v_w6981_v);
	assign v_w883_v = ~(v_w1775_v & v_w1772_v);
	assign v_w2507_v = ~(v_w992_v & v_w2429_v);
	assign v_w2188_v = ~(v_s218_v & v_w2187_v);
	assign v_w1125_v = ~(v_w1457_v | v_w1461_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s125_v<=0;
	end
	else
	begin
	v_s125_v<=v_w134_v;
	end
	end
	assign v_w5686_v = ~(v_s305_v & v_w528_v);
	assign v_w5040_v = ~(v_w5035_v | v_w5039_v);
	assign v_w6134_v = ~(v_w6132_v & v_w6133_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s15_v<=0;
	end
	else
	begin
	v_s15_v<=v_w16_v;
	end
	end
	assign v_w2129_v = ~(v_w2127_v & v_w2128_v);
	assign v_w2528_v = ~(v_w2526_v | v_w2527_v);
	assign v_w2548_v = ~(v_w2484_v & v_w2367_v);
	assign v_w5631_v = ~(v_w420_v & v_w2379_v);
	assign v_w7492_v = ~(v_w7326_v & v_w7491_v);
	assign v_w5947_v = ~(v_w5945_v | v_w5946_v);
	assign v_w6192_v = ~(v_w6191_v & v_w659_v);
	assign v_w830_v = ~(v_w982_v | v_w983_v);
	assign v_w2935_v = ~(v_w572_v);
	assign v_w2696_v = ~(v_w2694_v & v_w2695_v);
	assign v_w4974_v = ~(v_w4973_v & v_w673_v);
	assign v_w758_v = ~(v_w1777_v & v_w1785_v);
	assign v_w39_v = ~(v_w7134_v & v_w7135_v);
	assign v_w8126_v = v_w8125_v ^ v_keyinput_44_v;
	assign v_w4723_v = ~(v_w782_v | v_w4568_v);
	assign v_w3971_v = ~(v_w3767_v & v_w3970_v);
	assign v_w7890_v = ~(v_w651_v & v_w7777_v);
	assign v_w4380_v = ~(v_w4056_v & v_s392_v);
	assign v_w958_v = v_w956_v & v_w957_v;
	assign v_w782_v = ~(v_w781_v);
	assign v_w7759_v = ~(v_w7757_v & v_w7758_v);
	assign v_w7775_v = ~(v_w6795_v | v_w7774_v);
	assign v_w3318_v = ~(v_w3316_v & v_w3317_v);
	assign v_w5824_v = ~(v_w2117_v & v_w1064_v);
	assign v_w3420_v = ~(v_w3418_v | v_w3419_v);
	assign v_w3202_v = ~(v_w963_v & v_w2639_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s450_v<=0;
	end
	else
	begin
	v_s450_v<=v_w503_v;
	end
	end
	assign v_w4649_v = ~(v_w2448_v & v_w2706_v);
	assign v_w5351_v = ~(v_w4996_v | v_w5350_v);
	assign v_w7996_v = v_s464_v & v_s330_v;
	assign v_w2841_v = ~(v_w2840_v & v_w697_v);
	assign v_w2705_v = ~(v_w2355_v & v_s41_v);
	assign v_w1426_v = ~(v_w613_v & v_w1425_v);
	assign v_w3730_v = ~(v_w3618_v & v_w3729_v);
	assign v_w1109_v = ~(v_in8_v | v_w1201_v);
	assign v_w1221_v = ~(v_s103_v & v_w1103_v);
	assign v_w5404_v = ~(v_w1088_v | v_w2602_v);
	assign v_w6483_v = ~(v_w6481_v & v_w6482_v);
	assign v_w1576_v = ~(v_w8254_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s310_v<=0;
	end
	else
	begin
	v_s310_v<=v_w333_v;
	end
	end
	assign v_w4576_v = ~(v_w4575_v | v_w3629_v);
	assign v_w3738_v = ~(v_w1069_v | v_w3735_v);
	assign v_w4076_v = ~(v_w4074_v & v_w4075_v);
	assign v_w1903_v = ~(v_w1902_v & v_w962_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s21_v<=0;
	end
	else
	begin
	v_s21_v<=v_w23_v;
	end
	end
	assign v_w5421_v = ~(v_w2601_v & v_w968_v);
	assign v_w1225_v = ~(v_w612_v & v_s107_v);
	assign v_w5970_v = ~(v_w5968_v & v_w5969_v);
	assign v_w4732_v = ~(v_w674_v | v_w4731_v);
	assign v_w954_v = v_s111_v | v_s125_v;
	assign v_w562_v = v_w561_v;
	assign v_w6188_v = ~(v_w1514_v & v_w6160_v);
	assign v_w7809_v = ~(v_s415_v & v_w7742_v);
	assign v_w7014_v = ~(v_w6592_v & v_w1027_v);
	assign v_w5419_v = ~(v_w4822_v | v_w5123_v);
	assign v_w4833_v = ~(v_w4831_v & v_w4832_v);
	assign v_w1204_v = ~(v_w1202_v & v_w1203_v);
	assign v_w4083_v = ~(v_s256_v & v_w1037_v);
	assign v_w7255_v = ~(v_w680_v & v_w6585_v);
	assign v_w5922_v = ~(v_s340_v & v_w528_v);
	assign v_w1709_v = ~(v_w1707_v & v_w1708_v);
	assign v_w1276_v = ~(v_w1274_v & v_w1275_v);
	assign v_w6399_v = ~(v_w1440_v);
	assign v_w8089_v = v_w8088_v ^ v_keyinput_18_v;
	assign v_w4643_v = ~(v_w4642_v | v_w4528_v);
	assign v_w7187_v = ~(v_w1465_v | v_w529_v);
	assign v_w26_v = ~(v_w5676_v & v_w5677_v);
	assign v_w7613_v = ~(v_w7612_v | v_w1385_v);
	assign v_w1194_v = ~(v_w612_v & v_s29_v);
	assign v_w3193_v = ~(v_w3192_v & v_w697_v);
	assign v_w2831_v = ~(v_w2827_v);
	assign v_w5983_v = ~(v_w5979_v | v_w5982_v);
	assign v_w5748_v = ~(v_w5746_v & v_w5747_v);
	assign v_w1970_v = ~(v_w1966_v | v_w1969_v);
	assign v_w6764_v = ~(v_w6762_v & v_w6763_v);
	assign v_w2862_v = ~(v_w558_v & v_w2861_v);
	assign v_w5342_v = ~(v_w5340_v | v_w5341_v);
	assign v_w7309_v = v_w7305_v | v_w7308_v;
	assign v_w6417_v = v_s160_v ^ v_w6399_v;
	assign v_w5224_v = ~(v_w693_v | v_w2851_v);
	assign v_w7522_v = ~(v_w962_v | v_w680_v);
	assign v_w5727_v = ~(v_w5725_v & v_w5726_v);
	assign v_w2972_v = ~(v_w2970_v | v_w2971_v);
	assign v_w6334_v = ~(v_w6333_v & v_w6020_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s76_v<=0;
	end
	else
	begin
	v_s76_v<=v_w84_v;
	end
	end
	assign v_w5617_v = ~(v_w5555_v & v_w5546_v);
	assign v_w7902_v = ~(v_w651_v & v_w7814_v);
	assign v_w7376_v = ~(v_w680_v | v_w789_v);
	assign v_w3513_v = ~(v_w3508_v | v_w3512_v);
	assign v_w6332_v = v_w1644_v ^ v_w6331_v;
	assign v_w4000_v = ~(v_w3998_v & v_w3999_v);
	assign v_w5708_v = ~(v_w5707_v & v_w1280_v);
	assign v_w5833_v = ~(v_w2063_v & v_w2061_v);
	assign v_w6293_v = ~(v_w1610_v | v_w6271_v);
	assign v_w6317_v = v_w1644_v ^ v_w6316_v;
	assign v_w91_v = ~(v_w5598_v & v_w5599_v);
	assign v_w3608_v = ~(v_w3601_v | v_w3607_v);
	assign v_w4421_v = ~(v_w963_v | v_w4420_v);
	assign v_w3546_v = ~(v_w957_v & v_w3545_v);
	assign v_w7818_v = ~(v_w1065_v | v_w1782_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s311_v<=0;
	end
	else
	begin
	v_s311_v<=v_w334_v;
	end
	end
	assign v_w6185_v = ~(v_w6183_v ^ v_w6184_v);
	assign v_w652_v = ~(v_w2122_v & v_w2109_v);
	assign v_w6514_v = ~(v_w6510_v & v_w6513_v);
	assign v_w1244_v = ~(v_w612_v & v_s333_v);
	assign v_w3355_v = ~(v_w2956_v | v_w2620_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s357_v<=0;
	end
	else
	begin
	v_s357_v<=v_w395_v;
	end
	end
	assign v_w6378_v = ~(v_w6376_v & v_w6377_v);
	assign v_w1100_v = ~(v_w1498_v & v_w1499_v);
	assign v_w6540_v = ~(v_w6526_v & v_w6529_v);
	assign v_w4253_v = ~(v_w4252_v & v_w690_v);
	assign v_w6078_v = ~(v_w6047_v);
	assign v_w7412_v = ~(v_w687_v | v_w536_v);
	assign v_w801_v = ~(v_w1438_v & v_w1687_v);
	assign v_w6479_v = ~(v_w6474_v & v_w6478_v);
	assign v_w2629_v = ~(v_w2624_v);
	assign v_w6988_v = ~(v_w6979_v & v_w6987_v);
	assign v_w4127_v = ~(v_w2312_v & v_s241_v);
	assign v_w6272_v = ~(v_w1610_v ^ v_w6271_v);
	assign v_w2784_v = ~(v_w2782_v & v_w2783_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s463_v<=0;
	end
	else
	begin
	v_s463_v<=v_w516_v;
	end
	end
	assign v_w5396_v = ~(v_w4888_v & v_w5126_v);
	assign v_w1291_v = ~(v_w1290_v | v_w1180_v);
	assign v_w1745_v = ~(v_w1328_v | v_w1744_v);
	assign v_w542_v = ~(v_w540_v & v_w541_v);
	assign v_w5266_v = ~(v_w674_v & v_s430_v);
	assign v_w5115_v = ~(v_w5113_v | v_w5114_v);
	assign v_w2981_v = ~(v_w2980_v | v_w557_v);
	assign v_w3372_v = ~(v_w3063_v | v_w620_v);
	assign v_w4035_v = ~(v_w885_v | v_w4034_v);
	assign v_w5885_v = ~(v_w5693_v | v_w5884_v);
	assign v_w4496_v = ~(v_w4454_v & v_w4495_v);
	assign v_w785_v = ~(v_w1040_v & v_w1041_v);
	assign v_w8018_v = ~(v_w8002_v | v_w8017_v);
	assign v_w1529_v = ~(v_w666_v & v_s235_v);
	assign v_w8191_v = v_w5082_v & v_w5083_v;
	assign v_w3413_v = ~(v_w2588_v | v_w2620_v);
	assign v_w4122_v = ~(v_w690_v & v_w4121_v);
	assign v_w3366_v = ~(v_w2607_v & v_w2722_v);
	assign v_w3890_v = ~(v_w3888_v | v_w3889_v);
	assign v_w1069_v = ~(v_w1068_v);
	assign v_w4244_v = ~(v_s200_v ^ v_w2896_v);
	assign v_w7402_v = v_w7398_v | v_w7401_v;
	assign v_w3564_v = ~(v_w3560_v & v_w3563_v);
	assign v_w4261_v = ~(v_w4251_v | v_w4250_v);
	assign v_w4726_v = ~(v_w4725_v | v_w4589_v);
	assign v_w2666_v = ~(v_w2664_v & v_w2665_v);
	assign v_w1629_v = ~(v_w808_v | v_w1628_v);
	assign v_w4855_v = v_w2991_v ^ v_w4407_v;
	assign v_w3394_v = ~(v_w3392_v & v_w3393_v);
	assign v_w5647_v = ~(v_w420_v & v_w2890_v);
	assign v_w6772_v = ~(v_w6769_v & v_w6771_v);
	assign v_w3235_v = ~(v_w3233_v & v_w3234_v);
	assign v_w2488_v = v_w993_v | v_w2426_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s312_v<=0;
	end
	else
	begin
	v_s312_v<=v_w335_v;
	end
	end
	assign v_w1391_v = ~(v_s375_v ^ v_w1390_v);
	assign v_w1453_v = ~(v_w1451_v & v_w1452_v);
	assign v_w2735_v = ~(v_w2361_v | v_w2734_v);
	assign v_w3951_v = v_w3770_v | v_w3773_v;
	assign v_w1881_v = ~(v_w930_v & v_w1709_v);
	assign v_w6438_v = v_w1424_v | v_w6436_v;
	assign v_w4847_v = ~(v_w4845_v & v_w4846_v);
	assign v_w1085_v = ~(v_w2294_v | v_w1405_v);
	assign v_w6388_v = ~(v_s122_v ^ v_w6387_v);
	assign v_w979_v = ~(v_w766_v ^ v_w1101_v);
	assign v_w2246_v = ~(v_w2193_v | v_w604_v);
	assign v_w6326_v = ~(v_w1644_v ^ v_w6325_v);
	assign v_w5098_v = ~(v_w4863_v | v_w5097_v);
	assign v_w1505_v = ~(v_w613_v & v_w1504_v);
	assign v_w7538_v = ~(v_w687_v & v_w1803_v);
	assign v_w443_v = ~(v_w4760_v & v_w4775_v);
	assign v_w1648_v = ~(v_w1645_v | v_w1647_v);
	assign v_w183_v = ~(v_w5190_v & v_w5191_v);
	assign v_w590_v = ~(v_w972_v | v_w973_v);
	assign v_w7285_v = ~(v_w7283_v | v_w7284_v);
	assign v_w7049_v = ~(v_w7048_v & v_w758_v);
	assign v_w3878_v = ~(v_w3844_v | v_w3877_v);
	assign v_w6444_v = ~(v_w6442_v & v_w6443_v);
	assign v_w5508_v = ~(v_s187_v & v_w5386_v);
	assign v_w728_v = ~(v_w727_v | v_w643_v);
	assign v_w3777_v = ~(v_w3775_v | v_w3776_v);
	assign v_w6221_v = ~(v_w6214_v & v_w6220_v);
	assign v_w544_v = ~(v_s163_v ^ v_w543_v);
	assign v_w361_v = ~(v_w5642_v & v_w5643_v);
	assign v_w4178_v = ~(v_w4177_v & v_w692_v);
	assign v_w2335_v = ~(v_w2333_v | v_w2334_v);
	assign v_w3549_v = ~(v_w1083_v & v_w2993_v);
	assign v_w2856_v = ~(v_w2854_v | v_w2855_v);
	assign v_w5237_v = ~(v_w2571_v | v_w1_v);
	assign v_w4828_v = ~(v_w4456_v | v_w4557_v);
	assign v_w1706_v = ~(v_s393_v & v_w562_v);
	assign v_w8227_v = v_w8226_v ^ v_keyinput_111_v;
	assign v_w4674_v = ~(v_w2343_v & v_w4673_v);
	assign v_w8254_v = v_w8253_v ^ v_keyinput_127_v;
	assign v_w7901_v = ~(v_s31_v & v_w7876_v);
	assign v_w5838_v = ~(v_w1412_v | v_w2135_v);
	assign v_w4077_v = v_w4073_v ^ v_w4076_v;
	assign v_w1086_v = ~(v_w2958_v & v_w2962_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s360_v<=0;
	end
	else
	begin
	v_s360_v<=v_w399_v;
	end
	end
	assign v_w6630_v = ~(v_w6628_v | v_w6629_v);
	assign v_w4771_v = ~(v_w4769_v | v_w4770_v);
	assign v_w3595_v = ~(v_w3100_v & v_w3087_v);
	assign v_w2746_v = ~(v_w699_v & v_s179_v);
	assign v_w8072_v = v_w3866_v | v_w3867_v;
	assign v_w8023_v = ~(v_w8021_v | v_w8022_v);
	assign v_w6666_v = ~(v_w6663_v & v_w6665_v);
	assign v_w5219_v = ~(v_s346_v & v_w5140_v);
	assign v_w539_v = v_w604_v | v_w556_v;
	assign v_w831_v = ~(v_w830_v);
	assign v_w6111_v = ~(v_w1557_v | v_w6090_v);
	assign v_w616_v = ~(v_w605_v & v_w556_v);
	assign v_w7948_v = ~(v_w527_v & v_w1416_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s465_v<=0;
	end
	else
	begin
	v_s465_v<=v_w518_v;
	end
	end
	assign v_w4512_v = ~(v_w4510_v | v_w4511_v);
	assign v_w6594_v = ~(v_w655_v & v_w884_v);
	assign v_w3745_v = ~(v_w3743_v | v_w3744_v);
	assign v_w5063_v = ~(v_w2433_v);
	assign v_w1156_v = v_w1155_v | v_s339_v;
	assign v_w3998_v = ~(v_w3996_v | v_w3997_v);
	assign v_w7386_v = v_w7382_v | v_w7385_v;
	assign v_w3254_v = ~(v_s385_v & v_w1_v);
	assign v_w1445_v = ~(v_w1442_v | v_w1444_v);
	assign v_w2676_v = ~(v_w2674_v & v_w2675_v);
	assign v_w7727_v = ~(v_w1783_v & v_w1632_v);
	assign v_w7429_v = ~(v_w7402_v & v_w7428_v);
	assign v_w4262_v = ~(v_w4260_v | v_w4261_v);
	assign v_w948_v = ~(v_w648_v | v_w1844_v);
	assign v_w7805_v = ~(v_w7804_v | v_w6702_v);
	assign v_w440_v = ~(v_w4793_v & v_w4795_v);
	assign v_w4822_v = v_w4456_v ^ v_w4491_v;
	assign v_w8008_v = ~(v_w280_v | v_w8006_v);
	assign v_w5584_v = ~(v_s118_v & v_w676_v);
	assign v_w5488_v = ~(v_s422_v & v_w5386_v);
	assign v_w1060_v = ~(v_in6_v ^ v_w1195_v);
	assign v_w334_v = ~(v_w4180_v & v_w4186_v);
	assign v_w3517_v = ~(v_w3514_v & v_w3516_v);
	assign v_w6879_v = ~(v_w6877_v & v_w6878_v);
	assign v_w5531_v = v_w8225_v ^ v_keyinput_110_v;
	assign v_w6096_v = ~(v_s271_v & v_w1557_v);
	assign v_w1309_v = ~(v_w1307_v & v_w1308_v);
	assign v_w3007_v = ~(v_s105_v & v_w2355_v);
	assign v_w4725_v = v_w782_v ^ v_w4504_v;
	assign v_w2698_v = ~(v_w2478_v & v_w753_v);
	assign v_w1535_v = ~(v_w1051_v & v_s236_v);
	assign v_w2601_v = ~(v_w2257_v | v_w2235_v);
	assign v_w8209_v = v_w7810_v | v_w1919_v;
	assign v_w7958_v = ~(v_w527_v & v_w1362_v);
	assign v_w3621_v = v_w3620_v ^ v_w866_v;
	assign v_w5214_v = ~(v_w5212_v | v_w5213_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s381_v<=0;
	end
	else
	begin
	v_s381_v<=v_w427_v;
	end
	end
	assign v_w457_v = ~(v_w5797_v & v_w5804_v);
	assign v_w5324_v = ~(v_w5038_v & v_w5323_v);
	assign v_w1578_v = ~(v_s477_v & v_s7_v);
	assign v_w80_v = v_s72_v & v_w7107_v;
	assign v_w7565_v = ~(v_w1658_v & v_w1633_v);
	assign v_w6017_v = ~(v_w1190_v | v_w658_v);
	assign v_w5717_v = ~(v_w2056_v ^ v_w2057_v);
	assign v_w4386_v = ~(v_w4385_v & v_w692_v);
	assign v_w4543_v = ~(v_w3519_v & v_w4542_v);
	assign v_w1185_v = ~(v_w1181_v | v_w1184_v);
	assign v_w7604_v = v_w800_v & v_w1454_v;
	assign v_w4623_v = ~(v_w2342_v | v_w4622_v);
	assign v_w300_v = ~(v_w5048_v & v_w5053_v);
	assign v_w5988_v = ~(v_s440_v & v_w528_v);
	assign v_w2616_v = ~(v_w2612_v | v_w2615_v);
	assign v_w4286_v = ~(v_w2930_v & v_s352_v);
	assign v_w6846_v = ~(v_w6637_v | v_w6842_v);
	assign v_w6845_v = ~(v_w6838_v & v_w6844_v);
	assign v_w5262_v = ~(v_w5260_v | v_w5261_v);
	assign v_w1353_v = ~(v_w1352_v);
	assign v_w6981_v = ~(v_w1798_v & v_w1135_v);
	assign v_w3501_v = ~(v_w2401_v | v_w3500_v);
	assign v_w7935_v = ~(v_s325_v & v_w2143_v);
	assign v_w6007_v = ~(v_w2117_v & v_w1437_v);
	assign v_w3416_v = ~(v_w3121_v | v_w2562_v);
	assign v_w3824_v = ~(v_w2619_v | v_w3731_v);
	assign v_w5101_v = ~(v_w2447_v & v_w3216_v);
	assign v_w7321_v = ~(v_w7319_v | v_w7320_v);
	assign v_w6624_v = ~(v_w1787_v & v_w1297_v);
	assign v_w4483_v = ~(v_w3642_v | v_w4482_v);
	assign v_w4860_v = ~(v_w4858_v & v_w4859_v);
	assign v_w574_v = ~(v_w1573_v & v_w1574_v);
	assign v_w1388_v = v_w943_v & v_s7_v;
	assign v_w2758_v = ~(v_w1011_v | v_w617_v);
	assign v_w6174_v = ~(v_w6172_v & v_w6173_v);
	assign v_w3308_v = ~(v_w2639_v & v_w753_v);
	assign v_w7254_v = ~(v_w687_v & v_w7253_v);
	assign v_w6918_v = ~(v_w6641_v & v_w6917_v);
	assign v_w554_v = ~(v_w2238_v);
	assign v_w851_v = ~(v_w1014_v & v_w1015_v);
	assign v_w32_v = ~(v_w5674_v & v_w5675_v);
	assign v_w5834_v = ~(v_w5833_v ^ v_w628_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s224_v<=0;
	end
	else
	begin
	v_s224_v<=v_w237_v;
	end
	end
	assign v_w2741_v = v_w553_v ^ v_w2740_v;
	assign v_w5990_v = ~(v_w5988_v & v_w5989_v);
	assign v_w6956_v = ~(v_w6955_v & v_w1915_v);
	assign v_w1517_v = ~(v_w783_v ^ v_w542_v);
	assign v_w6873_v = ~(v_w758_v & v_w6872_v);
	assign v_w917_v = ~(v_w1115_v & v_w1116_v);
	assign v_w2107_v = ~(v_w2106_v);
	assign v_w6548_v = ~(v_w6546_v | v_w6547_v);
	assign v_w70_v = v_s62_v & v_w7107_v;
	assign v_w2606_v = ~(v_w2605_v & v_w1037_v);
	assign v_w3640_v = ~(v_w3639_v);
	assign v_w5276_v = ~(v_w3678_v ^ v_w5275_v);
	assign v_w3230_v = ~(v_w3228_v | v_w3229_v);
	assign v_w2364_v = ~(v_w2361_v | v_w2363_v);
	assign v_w3247_v = v_w3243_v ^ v_w3246_v;
	assign v_w1680_v = ~(v_w1663_v & v_w1679_v);
	assign v_w2436_v = ~(v_w2435_v & v_w2407_v);
	assign v_w362_v = ~(v_w7193_v & v_w7194_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s391_v<=0;
	end
	else
	begin
	v_s391_v<=v_w440_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s519_v<=0;
	end
	else
	begin
	v_s519_v<=v_w528_v;
	end
	end
	assign v_w4919_v = ~(v_w2261_v | v_w2906_v);
	assign v_w4631_v = ~(v_w3095_v | v_w2370_v);
	assign v_w5946_v = ~(v_w1125_v | v_w2138_v);
	assign v_w7709_v = ~(v_w7707_v | v_w7708_v);
	assign v_w3337_v = ~(v_w1139_v & v_w3336_v);
	assign v_w423_v = ~(v_w3294_v & v_w3296_v);
	assign v_w1016_v = ~(v_w1011_v);
	assign v_w3556_v = ~(v_w2753_v & v_w1016_v);
	assign v_w6672_v = ~(v_w6671_v & v_w655_v);
	assign v_w1262_v = ~(v_w1260_v & v_w1261_v);
	assign v_w679_v = v_w687_v;
	assign v_w4677_v = ~(v_w4675_v & v_w4676_v);
	assign v_w1682_v = ~(v_w1681_v & v_w901_v);
	assign v_w4126_v = v_w4116_v ^ v_s239_v;
	assign v_w3764_v = ~(v_w852_v & v_w3732_v);
	assign v_w2602_v = ~(v_w2601_v);
	assign v_w8144_v = ~(v_w2663_v | v_w2672_v);
	assign v_w4920_v = ~(v_w4918_v | v_w4919_v);
	assign v_w157_v = v_s148_v & v_w5134_v;
	assign v_w7676_v = ~(v_w8190_v);
	assign v_w1775_v = ~(v_w1774_v);
	assign v_w6792_v = ~(v_w1373_v | v_w1797_v);
	assign v_w3710_v = ~(v_w3708_v | v_w3709_v);
	assign v_w2314_v = ~(v_w568_v | v_w2313_v);
	assign v_w1663_v = ~(v_w1472_v & v_w1662_v);
	assign v_w6914_v = ~(v_w6913_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s110_v<=0;
	end
	else
	begin
	v_s110_v<=v_w118_v;
	end
	end
	assign v_w891_v = ~(v_w716_v & v_s7_v);
	assign v_w5739_v = ~(v_w892_v & v_w1632_v);
	assign v_w4794_v = v_w1079_v ^ v_w4410_v;
	assign v_w4263_v = v_w4259_v ^ v_w4262_v;
	assign v_w5764_v = ~(v_w5762_v & v_w5763_v);
	assign v_w4008_v = ~(v_w3749_v & v_w4007_v);
	assign v_w7195_v = ~(v_w1626_v | v_w528_v);
	assign v_w2728_v = ~(v_w2726_v & v_w2727_v);
	assign v_w1250_v = ~(v_s208_v & v_w1103_v);
	assign v_w5612_v = ~(v_s23_v & v_w676_v);
	assign v_w261_v = ~(v_w7919_v & v_w7920_v);
	assign v_w5802_v = ~(v_w5800_v & v_w5801_v);
	assign v_w3816_v = ~(v_w2827_v & v_w3732_v);
	assign v_w1395_v = ~(v_w666_v & v_s108_v);
	assign v_w4808_v = ~(v_w4797_v & v_w4807_v);
	assign v_w2584_v = ~(v_w699_v & v_s220_v);
	assign v_w4622_v = v_w4616_v ^ v_w4418_v;
	assign v_w1338_v = ~(v_w918_v & v_w1337_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s425_v<=0;
	end
	else
	begin
	v_s425_v<=v_w476_v;
	end
	end
	assign v_w1743_v = ~(v_w1738_v & v_w1742_v);
	assign v_w2282_v = ~(v_w2275_v & v_w2281_v);
	assign v_w5476_v = ~(v_w4705_v | v_w5123_v);
	assign v_w5274_v = ~(v_w3118_v | v_w963_v);
	assign v_w7513_v = ~(v_w1337_v | v_w7505_v);
	assign v_w5721_v = ~(v_w1446_v | v_w2135_v);
	assign v_w2422_v = ~(v_w2420_v & v_w2421_v);
	assign v_w4916_v = ~(v_w674_v & v_s331_v);
	assign v_w6331_v = ~(v_w6329_v & v_w6330_v);
	assign v_w3651_v = ~(v_w2461_v & v_w2427_v);
	assign v_w1843_v = ~(v_w1548_v & v_w1842_v);
	assign v_w4477_v = ~(v_w3639_v | v_w4476_v);
	assign v_w1255_v = ~(v_w1253_v & v_w1254_v);
	assign v_w8077_v = ~(v_w7460_v | v_w7461_v);
	assign v_w4977_v = ~(v_w4976_v & v_w878_v);
	assign v_w4469_v = ~(v_w4459_v & v_w4468_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s239_v<=0;
	end
	else
	begin
	v_s239_v<=v_w252_v;
	end
	end
	assign v_w3398_v = ~(v_w3396_v & v_w3397_v);
	assign v_w6861_v = ~(v_w6856_v & v_w6860_v);
	assign v_w7200_v = ~(v_w1607_v | v_w7117_v);
	assign v_w206_v = ~(v_w5644_v & v_w5645_v);
	assign v_w1860_v = ~(v_w726_v | v_w1859_v);
	assign v_w2304_v = ~(v_s276_v | v_w2288_v);
	assign v_w3572_v = ~(v_w3564_v & v_w3571_v);
	assign v_w6902_v = ~(v_w1642_v | v_w6608_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s441_v<=0;
	end
	else
	begin
	v_s441_v<=v_w493_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s333_v<=0;
	end
	else
	begin
	v_s333_v<=v_w361_v;
	end
	end
	assign v_w4657_v = ~(v_w4656_v & v_w878_v);
	assign v_w1479_v = ~(v_s213_v & v_w562_v);
	assign v_w3889_v = ~(v_w3885_v | v_w3882_v);
	assign v_w3452_v = ~(v_w3451_v);
	assign v_w6898_v = ~(v_w6638_v | v_w6894_v);
	assign v_w844_v = v_w843_v & v_s476_v;
	assign v_w1959_v = ~(v_w1957_v & v_w1958_v);
	assign v_w6611_v = ~(v_s449_v & v_w656_v);
	assign v_w2055_v = ~(v_w2010_v | v_w631_v);
	assign v_w3241_v = ~(v_w3239_v & v_w3240_v);
	assign v_w624_v = ~(v_w3023_v | v_w3027_v);
	assign v_w4460_v = ~(v_w2382_v | v_w2474_v);
	assign v_w4355_v = ~(v_w4330_v & v_w4333_v);
	assign v_w7974_v = ~(v_w527_v & v_w1762_v);
	assign v_w5513_v = ~(v_w5511_v | v_w5512_v);
	assign v_w2506_v = ~(v_w558_v & v_w2417_v);
	assign v_w2493_v = ~(v_w2426_v | v_w538_v);
	assign v_w6246_v = ~(v_w6245_v & v_w659_v);
	assign v_w2091_v = ~(v_w8104_v);
	assign v_w7789_v = ~(v_w6754_v & v_w7788_v);
	assign v_w3826_v = ~(v_w2619_v | v_w3735_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s1_v<=0;
	end
	else
	begin
	v_s1_v<=v_w1_v;
	end
	end
	assign v_w753_v = ~(v_w860_v & v_w861_v);
	assign v_w7951_v = ~(v_s103_v & v_w2143_v);
	assign v_w235_v = ~(v_w5634_v & v_w5635_v);
	assign v_w1155_v = v_s337_v | v_w1154_v;
	assign v_w4885_v = v_w1017_v ^ v_w4405_v;
	assign v_w6948_v = ~(v_w6947_v);
	assign v_w3771_v = ~(v_w761_v & v_w3732_v);
	assign v_w2815_v = v_s313_v ^ v_w2641_v;
	assign v_w5359_v = ~(v_w5357_v & v_w5358_v);
	assign v_w6896_v = ~(v_w1862_v ^ v_w1661_v);
	assign v_w8245_v = v_w8244_v ^ v_keyinput_122_v;
	assign v_w5183_v = ~(v_w1354_v & v_w5146_v);
	assign v_w4851_v = ~(v_w4844_v & v_w4850_v);
	assign v_w4969_v = ~(v_w2448_v & v_w2618_v);
	assign v_w2757_v = ~(v_w2756_v & v_w569_v);
	assign v_w3526_v = ~(v_w2819_v | v_w2831_v);
	assign v_w7462_v = ~(v_w8078_v);
	assign v_w2448_v = v_w2447_v;
	assign v_w5863_v = ~(v_w1397_v | v_w2135_v);
	assign v_w8041_v = ~(v_w7989_v | v_w8040_v);
	assign v_w6513_v = ~(v_w6511_v & v_w6512_v);
	assign v_w7997_v = ~(v_s463_v | v_s317_v);
	assign v_w1104_v = v_w1103_v & v_in33_v;
	assign v_w113_v = ~(v_w5592_v & v_w5593_v);
	assign v_w693_v = ~(v_s1_v);
	assign v_w7060_v = ~(v_s272_v | v_w6571_v);
	assign v_w1411_v = ~(v_w1409_v & v_w1410_v);
	assign v_w7705_v = ~(v_s225_v & v_w7667_v);
	assign v_w7207_v = ~(v_w1490_v | v_w528_v);
	assign v_w575_v = ~(v_w573_v | v_w574_v);
	assign v_o13_v = ~(v_w8024_v ^ v_w8025_v);
	assign v_w3550_v = ~(v_w3548_v & v_w3549_v);
	assign v_w174_v = ~(v_w5170_v & v_w5171_v);
	assign v_w4728_v = ~(v_w2448_v & v_w2738_v);
	assign v_w33_v = ~(v_w7130_v & v_w7131_v);
	assign v_w3453_v = ~(v_s6_v & v_w612_v);
	assign v_w1474_v = ~(v_s302_v ^ v_w1473_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s453_v<=0;
	end
	else
	begin
	v_s453_v<=v_w506_v;
	end
	end
	assign v_w6716_v = ~(v_w6712_v & v_w6715_v);
	assign v_w3168_v = ~(v_w3125_v | v_w3167_v);
	assign v_w5622_v = ~(v_s264_v & v_w695_v);
	assign v_w3854_v = ~(v_w2326_v & v_w3732_v);
	assign v_w1753_v = ~(v_w8184_v);
	assign v_w2509_v = ~(v_w2505_v | v_w2508_v);
	assign v_w6160_v = ~(v_w6158_v & v_w6159_v);
	assign v_w5976_v = ~(v_w5975_v & v_w2113_v);
	assign v_w4616_v = ~(v_w871_v);
	assign v_w7344_v = ~(v_w7342_v | v_w7343_v);
	assign v_w6314_v = ~(v_s205_v & v_w1626_v);
	assign v_w5697_v = ~(v_w5695_v | v_w5696_v);
	assign v_w8102_v = v_in6_v | v_w1195_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s335_v<=0;
	end
	else
	begin
	v_s335_v<=v_w364_v;
	end
	end
	assign v_w1497_v = ~(v_w1180_v | v_w1496_v);
	assign v_w7575_v = ~(v_w6824_v & v_w7574_v);
	assign v_w1620_v = ~(v_w1618_v & v_w1619_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s57_v<=0;
	end
	else
	begin
	v_s57_v<=v_w65_v;
	end
	end
	assign v_w7437_v = ~(v_w7435_v | v_w7436_v);
	assign v_w2368_v = ~(v_w2367_v);
	assign v_w3940_v = ~(v_w3936_v | v_w3939_v);
	assign v_w7044_v = ~(v_w7043_v & v_w655_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s200_v<=0;
	end
	else
	begin
	v_s200_v<=v_w213_v;
	end
	end
	assign v_w5334_v = ~(v_w5332_v & v_w5333_v);
	assign v_w6496_v = ~(v_s406_v & v_w6457_v);
	assign v_w7390_v = ~(v_w7388_v | v_w7389_v);
	assign v_w1408_v = ~(v_w613_v & v_w1407_v);
	assign v_w2826_v = ~(v_w1607_v | v_w2294_v);
	assign v_w6009_v = ~(v_w1428_v | v_w2135_v);
	assign v_w3910_v = ~(v_w3808_v & v_w3909_v);
	assign v_w4383_v = ~(v_w4381_v | v_w4382_v);
	assign v_w766_v = ~(v_w765_v);
	assign v_w5674_v = ~(v_s29_v & v_w695_v);
	assign v_w291_v = ~(v_w7061_v & v_w7062_v);
	assign v_w2051_v = ~(v_w2049_v & v_w2050_v);
	assign v_w4193_v = ~(v_w4192_v & v_w692_v);
	assign v_w1985_v = ~(v_w1983_v & v_w1984_v);
	assign v_w5602_v = ~(v_s42_v & v_w676_v);
	assign v_w2570_v = ~(v_w2294_v | v_w1488_v);
	assign v_w6069_v = ~(v_s270_v & v_w528_v);
	assign v_w6423_v = ~(v_w5712_v | v_w6422_v);
	assign v_w4665_v = ~(v_w674_v & v_s421_v);
	assign v_w1364_v = ~(v_w1119_v & v_w1363_v);
	assign v_w350_v = ~(v_w6942_v & v_w6943_v);
	assign v_w207_v = ~(v_w7741_v & v_w7743_v);
	assign v_w2462_v = ~(v_w2335_v | v_w2426_v);
	assign v_w5792_v = ~(v_w5791_v & v_w5703_v);
	assign v_w6714_v = ~(v_w6713_v);
	assign v_w1021_v = ~(v_w1020_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s180_v<=0;
	end
	else
	begin
	v_s180_v<=v_w193_v;
	end
	end
	assign v_w6638_v = ~(v_w8188_v);
	assign v_w4290_v = ~(v_w692_v & v_w4289_v);
	assign v_w1424_v = ~(v_s368_v ^ v_w1423_v);
	assign v_w877_v = ~(v_w554_v & v_w2233_v);
	assign v_w180_v = ~(v_w5178_v & v_w5179_v);
	assign v_w5884_v = ~(v_w5883_v ^ v_w611_v);
	assign v_w379_v = ~(v_w6893_v & v_w6905_v);
	assign v_w4016_v = ~(v_w4015_v & v_w881_v);
	assign v_w1550_v = ~(v_w1051_v & v_s246_v);
	assign v_w2708_v = ~(v_w2698_v & v_w2707_v);
	assign v_w2523_v = ~(v_w2482_v ^ v_w2486_v);
	assign v_w1836_v = ~(v_w1834_v | v_w1835_v);
	assign v_w7845_v = ~(v_w6570_v & v_w7844_v);
	assign v_w5837_v = ~(v_w5835_v & v_w5836_v);
	assign v_w54_v = v_s46_v & v_w7107_v;
	assign v_w6825_v = v_w6824_v ^ v_w1876_v;
	assign v_w45_v = ~(v_w7961_v & v_w7962_v);
	assign v_w7418_v = v_w7414_v | v_w7417_v;
	assign v_w2277_v = ~(v_w2276_v & v_w2170_v);
	assign v_w6268_v = ~(v_w6266_v | v_w6267_v);
	assign v_w4515_v = ~(v_w1008_v | v_w4514_v);
	assign v_w1827_v = ~(v_w1101_v | v_w765_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s185_v<=0;
	end
	else
	begin
	v_s185_v<=v_w198_v;
	end
	end
	assign v_w1366_v = ~(v_w874_v & v_s402_v);
	assign v_w220_v = ~(v_w7870_v & v_w7871_v);
	assign v_w2284_v = ~(v_w1037_v);
	assign v_w1015_v = ~(v_w2300_v & v_w1339_v);
	assign v_w7208_v = ~(v_w7117_v | v_w1488_v);
	assign v_w7971_v = ~(v_s14_v & v_w2143_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s506_v<=0;
	end
	else
	begin
	v_s506_v<=v_w376_v;
	end
	end
	assign v_w5234_v = ~(v_w5232_v | v_w5233_v);
	assign v_w6779_v = ~(v_w1883_v | v_w6579_v);
	assign v_w4807_v = ~(v_w4804_v | v_w4806_v);
	assign v_w5540_v = ~(v_w5286_v & v_w5539_v);
	assign v_w3392_v = ~(v_w2327_v & v_w2639_v);
	assign v_w2905_v = ~(v_w2903_v & v_w2904_v);
	assign v_w7076_v = ~(v_w1798_v & v_w578_v);
	assign v_w902_v = ~(v_w900_v & v_w901_v);
	assign v_w6040_v = ~(v_w6032_v | v_w6039_v);
	assign v_w3062_v = ~(v_w3052_v & v_w3061_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s268_v<=0;
	end
	else
	begin
	v_s268_v<=v_w285_v;
	end
	end
	assign v_w3020_v = ~(v_w864_v | v_w616_v);
	assign v_w1565_v = ~(v_s35_v & v_w670_v);
	assign v_w1942_v = ~(v_s56_v | v_s55_v);
	assign v_w3724_v = ~(v_w3723_v & v_w3613_v);
	assign v_w1577_v = ~(v_s264_v & v_w614_v);
	assign v_w688_v = ~(v_w1136_v & v_w1037_v);
	assign v_w4800_v = ~(v_w4560_v & v_w878_v);
	assign v_w2034_v = v_w2031_v & v_w2033_v;
	assign v_w899_v = v_w897_v & v_w898_v;
	assign v_w179_v = ~(v_w5182_v & v_w5183_v);
	assign v_w1848_v = ~(v_w1845_v & v_w1847_v);
	assign v_w2853_v = ~(v_w2852_v & v_w569_v);
	assign v_w3884_v = ~(v_w3735_v | v_w2585_v);
	assign v_w6387_v = v_w1667_v ^ v_w6386_v;
	assign v_w3968_v = ~(v_w3966_v & v_w3967_v);
	assign v_w6464_v = v_w6457_v ^ v_w6463_v;
	assign v_w7598_v = ~(v_w8234_v);
	assign v_w4334_v = v_w4330_v ^ v_w4333_v;
	assign v_w6583_v = ~(v_w3477_v & v_w809_v);
	assign v_w5278_v = ~(v_w5272_v & v_w5277_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s172_v<=0;
	end
	else
	begin
	v_s172_v<=v_w184_v;
	end
	end
	assign v_w5634_v = ~(v_s222_v & v_w695_v);
	assign v_w4535_v = ~(v_w3641_v);
	assign v_w467_v = ~(v_w7815_v & v_w7816_v);
	assign v_w5667_v = ~(v_w4082_v & v_w3077_v);
	assign v_w7363_v = ~(v_w7361_v | v_w7362_v);
	assign v_w5664_v = ~(v_s78_v & v_w695_v);
	assign v_w213_v = ~(v_w5578_v & v_w5579_v);
	assign v_w5953_v = ~(v_w5949_v | v_w5952_v);
	assign v_w7409_v = ~(v_w7407_v | v_w7408_v);
	assign v_w4369_v = ~(v_w3403_v | v_w4368_v);
	assign v_w2184_v = ~(v_w2180_v & v_w2183_v);
	assign v_w7881_v = ~(v_s160_v & v_w7876_v);
	assign v_w8052_v = ~(v_w547_v & v_w559_v);
	assign v_w7824_v = ~(v_w6652_v | v_w7823_v);
	assign v_w5036_v = v_w2309_v ^ v_w2338_v;
	assign v_w3173_v = ~(v_w3172_v | v_w2620_v);
	assign v_w6172_v = ~(v_w1514_v & v_w6171_v);
	assign v_w3014_v = ~(v_s103_v & v_w564_v);
	assign v_w678_v = v_w677_v | v_w8_v;
	assign v_w5221_v = ~(v_w2897_v | v_w1_v);
	assign v_w7587_v = ~(v_w1063_v & v_w7586_v);
	assign v_w1289_v = ~(v_w806_v ^ v_w807_v);
	assign v_w6613_v = ~(v_w6611_v & v_w6612_v);
	assign v_w6275_v = ~(v_s215_v & v_w1474_v);
	assign v_w7338_v = ~(v_w687_v | v_w1453_v);
	assign v_w3373_v = v_w3372_v ^ v_w3066_v;
	assign v_w4927_v = ~(v_w4926_v | v_w4589_v);
	assign v_w3999_v = ~(v_w3735_v & v_w2671_v);
	assign v_w2786_v = ~(v_w565_v & v_s90_v);
	assign v_w3831_v = ~(v_w2297_v & v_w3731_v);
	assign v_w378_v = ~(v_w5856_v & v_w5864_v);
	assign v_w2377_v = ~(v_w2375_v & v_w2376_v);
	assign v_w5517_v = ~(v_w4863_v | v_w4599_v);
	assign v_w1008_v = ~(v_w1006_v | v_w1007_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s70_v<=0;
	end
	else
	begin
	v_s70_v<=v_w78_v;
	end
	end
	assign v_w5975_v = ~(v_w599_v ^ v_w2065_v);
	assign v_w2814_v = ~(v_w2812_v & v_w2813_v);
	assign v_w3627_v = ~(v_w3626_v);
	assign v_w4497_v = ~(v_w4453_v | v_w4496_v);
	assign v_w2680_v = v_w2679_v ^ v_w553_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s66_v<=0;
	end
	else
	begin
	v_s66_v<=v_w74_v;
	end
	end
	assign v_w2986_v = ~(v_w2985_v & v_w569_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s502_v<=0;
	end
	else
	begin
	v_s502_v<=v_w362_v;
	end
	end
	assign v_w6965_v = ~(v_w1856_v | v_w1797_v);
	assign v_w1768_v = ~(v_w809_v & v_w1767_v);
	assign v_w763_v = ~(v_w3081_v | v_w817_v);
	assign v_w1732_v = ~(v_w1727_v | v_w1731_v);
	assign v_w2140_v = ~(v_s448_v & v_w529_v);
	assign v_w5719_v = ~(v_w892_v & v_w1681_v);
	assign v_w5472_v = ~(v_s184_v & v_w5386_v);
	assign v_w275_v = ~(v_w4053_v & v_w4055_v);
	assign v_w6065_v = ~(v_w6029_v | v_w6064_v);
	assign v_w5364_v = ~(v_w2601_v & v_w2831_v);
	assign v_w4839_v = ~(v_w2976_v & v_w2347_v);
	assign v_w6788_v = ~(v_w6787_v & v_w884_v);
	assign v_o16_v = ~(v_w8015_v ^ v_w8016_v);
	assign v_w4086_v = ~(v_w4082_v & v_w4085_v);
	assign v_w4917_v = ~(v_w2265_v & v_w2901_v);
	assign v_w2691_v = ~(v_w558_v & v_w2690_v);
	assign v_w1669_v = ~(v_w1668_v & v_w613_v);
	assign v_w4475_v = ~(v_w2863_v | v_w2861_v);
	assign v_w6402_v = ~(v_w6401_v & v_w6020_v);
	assign v_w1197_v = ~(v_w612_v & v_s34_v);
	assign v_w3432_v = ~(v_w871_v & v_w2639_v);
	assign v_w2382_v = ~(v_w2380_v | v_w2381_v);
	assign v_w1955_v = ~(v_w1947_v & v_w1954_v);
	assign v_w4758_v = ~(v_w4756_v & v_w4757_v);
	assign v_w4404_v = ~(v_w2916_v & v_w4403_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s284_v<=0;
	end
	else
	begin
	v_s284_v<=v_w303_v;
	end
	end
	assign v_w5139_v = ~(v_w1_v & v_w3467_v);
	assign v_w7713_v = ~(v_w7693_v | v_w6969_v);
	assign v_w3892_v = ~(v_w3828_v & v_w3825_v);
	assign v_w3655_v = ~(v_w2441_v & v_w3654_v);
	assign v_w1441_v = ~(v_w613_v & v_w1440_v);
	assign v_w3819_v = ~(v_w3735_v & v_w2833_v);
	assign v_w3897_v = ~(v_w3815_v & v_w3896_v);
	assign v_w4523_v = ~(v_w4521_v | v_w4522_v);
	assign v_w1563_v = ~(v_w1062_v ^ v_s157_v);
	assign v_w4589_v = ~(v_w4588_v);
	assign v_w4522_v = ~(v_w3100_v | v_w3098_v);
	assign v_w4063_v = ~(v_w4062_v & v_w692_v);
	assign v_w2639_v = ~(v_w2261_v & v_w2638_v);
	assign v_w5747_v = ~(v_w2137_v & v_w944_v);
	assign v_w6952_v = ~(v_w1787_v & v_w1135_v);
	assign v_w5073_v = ~(v_w5061_v & v_w5072_v);
	assign v_w5656_v = ~(v_s393_v & v_w695_v);
	assign v_w4559_v = ~(v_w3553_v & v_w4558_v);
	assign v_w4705_v = v_w4507_v ^ v_w3631_v;
	assign v_w7942_v = ~(v_w527_v & v_w1678_v);
	assign v_w317_v = ~(v_w4144_v & v_w4150_v);
	assign v_w6625_v = v_w934_v ^ v_w1906_v;
	assign v_w1067_v = ~(v_w1066_v);
	assign v_w1708_v = ~(v_w1075_v & v_w895_v);
	assign v_w7364_v = v_w7360_v | v_w7363_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s228_v<=0;
	end
	else
	begin
	v_s228_v<=v_w241_v;
	end
	end
	assign v_w1439_v = ~(v_s366_v & v_w562_v);
	assign v_w1944_v = ~(v_s60_v | v_s62_v);
	assign v_w5875_v = ~(v_w5873_v | v_w5874_v);
	assign v_w6469_v = ~(v_w1424_v & v_w6428_v);
	assign v_w7387_v = ~(v_w7382_v & v_w7385_v);
	assign v_w2614_v = ~(v_w337_v ^ v_w2613_v);
	assign v_w292_v = ~(v_w7921_v & v_w7922_v);
	assign v_w1842_v = ~(v_w1832_v & v_w1841_v);
	assign v_w1266_v = ~(v_s237_v & v_w1192_v);
	assign v_w1271_v = ~(v_w1269_v & v_w1270_v);
	assign v_w403_v = ~(v_w3268_v & v_w3274_v);
	assign v_w5705_v = ~(v_w2096_v | v_w2098_v);
	assign v_w4341_v = ~(v_w4337_v & v_w4340_v);
	assign v_w3696_v = ~(v_w3504_v | v_w2444_v);
	assign v_w2369_v = ~(v_w1037_v | v_w2242_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s422_v<=0;
	end
	else
	begin
	v_s422_v<=v_w473_v;
	end
	end
	assign v_w7648_v = ~(v_s12_v & v_w7647_v);
	assign v_w1961_v = ~(v_w1956_v & v_w1960_v);
	assign v_w7542_v = ~(v_w7534_v | v_w7541_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s303_v<=0;
	end
	else
	begin
	v_s303_v<=v_w326_v;
	end
	end
	assign v_w4824_v = ~(v_w4821_v | v_w4823_v);
	assign v_w5157_v = v_w5140_v & v_s18_v;
	assign v_w4901_v = ~(v_w2347_v & v_w2922_v);
	assign v_w2727_v = ~(v_w2484_v & v_w2722_v);
	assign v_w6681_v = ~(v_w758_v & v_w6679_v);
	assign v_w472_v = ~(v_w4672_v & v_w4674_v);
	assign v_w6863_v = ~(v_w6861_v | v_w6862_v);
	assign v_w2020_v = ~(v_w1837_v | v_w723_v);
	assign v_w40_v = ~(v_s483_v);
	assign v_w5881_v = ~(v_w5879_v & v_w5880_v);
	assign v_w1573_v = ~(v_s86_v & v_w670_v);
	assign v_w545_v = ~(v_w732_v & v_w733_v);
	assign v_w13_v = ~(v_w7651_v | v_w7652_v);
	assign v_w2366_v = ~(v_w699_v & v_s228_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s3_v<=0;
	end
	else
	begin
	v_s3_v<=v_w3_v;
	end
	end
	assign v_w841_v = ~(v_w769_v | v_w1042_v);
	assign v_w4372_v = ~(v_w2756_v | v_s389_v);
	assign v_w1452_v = ~(v_w875_v & v_s341_v);
	assign v_w5641_v = ~(v_w420_v & v_w2863_v);
	assign v_w907_v = ~(v_s388_v & v_w693_v);
	assign v_w5923_v = ~(v_w662_v & v_w1126_v);
	assign v_w6463_v = ~(v_w6461_v & v_w6462_v);
	assign v_w3396_v = ~(v_w1139_v & v_w3395_v);
	assign v_w3757_v = ~(v_w754_v & v_w3732_v);
	assign v_w6236_v = ~(v_s306_v & v_w6218_v);
	assign v_w6095_v = ~(v_w6093_v | v_w6094_v);
	assign v_w4217_v = v_w4213_v ^ v_w4216_v;
	assign v_w1339_v = ~(v_w1055_v ^ v_w1056_v);
	assign v_w3844_v = ~(v_w3836_v & v_w3843_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s328_v<=0;
	end
	else
	begin
	v_s328_v<=v_w356_v;
	end
	end
	assign v_w5417_v = ~(v_w683_v & v_w5416_v);
	assign v_w3729_v = ~(v_w2454_v | v_w3728_v);
	assign v_w4147_v = ~(v_w4117_v & v_w4120_v);
	assign v_w4196_v = ~(v_w4193_v & v_w4195_v);
	assign v_w2535_v = ~(v_w2529_v | v_w2532_v);
	assign v_w5683_v = ~(v_w4082_v & v_w3451_v);
	assign v_w8247_v = v_w2261_v | v_w2702_v;
	assign v_w5897_v = ~(v_w2044_v & v_w5896_v);
	assign v_w7233_v = ~(v_w7231_v | v_w7232_v);
	assign v_w2300_v = ~(v_w2294_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s174_v<=0;
	end
	else
	begin
	v_s174_v<=v_w187_v;
	end
	end
	assign v_w181_v = ~(v_s488_v);
	assign v_w2950_v = ~(v_w2355_v & v_s118_v);
	assign v_w6296_v = ~(v_s205_v & v_w888_v);
	assign v_w852_v = ~(v_w851_v);
	assign v_w4527_v = ~(v_w4526_v | v_w674_v);
	assign v_w4586_v = ~(v_w2448_v & v_w3100_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s225_v<=0;
	end
	else
	begin
	v_s225_v<=v_w238_v;
	end
	end
	assign v_w1396_v = ~(v_w1394_v & v_w1395_v);
	assign v_w846_v = ~(v_w1387_v & v_w1393_v);
	assign v_w1429_v = ~(v_w1428_v | v_w1180_v);
	assign v_w996_v = ~(v_w994_v & v_w995_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s493_v<=0;
	end
	else
	begin
	v_s493_v<=v_w279_v;
	end
	end
	assign v_w4444_v = ~(v_w674_v | v_w2370_v);
	assign v_w2745_v = ~(v_w2741_v | v_w2744_v);
	assign v_w7350_v = ~(v_w687_v | v_w1096_v);
	assign v_w7722_v = ~(v_w6959_v & v_w7721_v);
	assign v_w5780_v = ~(v_w5707_v & v_w1484_v);
	assign v_w4926_v = v_w4476_v ^ v_w3639_v;
	assign v_w3927_v = ~(v_w3784_v & v_w3926_v);
	assign v_w1850_v = ~(v_w1829_v & v_w1849_v);
	assign v_w3508_v = ~(v_w3507_v);
	assign v_w3713_v = ~(v_w3712_v & v_w3563_v);
	assign v_w4403_v = ~(v_w2861_v | v_w4402_v);
	assign v_w3618_v = ~(v_w3452_v & v_w3469_v);
	assign v_w5848_v = ~(v_w5847_v ^ v_w646_v);
	assign v_w6777_v = ~(v_w6775_v | v_w6776_v);
	assign v_w5941_v = ~(v_w5935_v & v_w5940_v);
	assign v_w6960_v = ~(v_w656_v | v_w6959_v);
	assign v_w5855_v = ~(v_w1418_v | v_w5734_v);
	assign v_w3949_v = ~(v_w3947_v & v_w3948_v);
	assign v_w1270_v = ~(v_w612_v & v_s242_v);
	assign v_w6882_v = ~(v_w6880_v & v_w6881_v);
	assign v_w4471_v = ~(v_w3645_v | v_w4470_v);
	assign v_w5310_v = ~(v_w4863_v | v_w5092_v);
	assign v_w3136_v = ~(v_w2952_v & v_w2634_v);
	assign v_w2700_v = ~(v_w2358_v & v_s421_v);
	assign v_w3071_v = ~(v_w2358_v & v_s410_v);
	assign v_w4113_v = ~(v_w690_v & v_w4112_v);
	assign v_w7960_v = ~(v_w527_v & v_w1350_v);
	assign v_w8096_v = v_w8095_v ^ v_keyinput_23_v;
	assign v_w8070_v = ~(v_w3492_v | v_w3542_v);
	assign v_w1456_v = ~(v_w875_v & v_s344_v);
	assign v_w6955_v = ~(v_w6909_v ^ v_w923_v);
	assign v_w3446_v = ~(v_w3442_v | v_w3445_v);
	assign v_w8235_v = ~(v_w1259_v & v_w739_v);
	assign v_w6549_v = ~(v_w1701_v & v_w6515_v);
	assign v_w4389_v = ~(v_w3018_v & v_s391_v);
	assign v_w5066_v = ~(v_w5065_v & v_w878_v);
	assign v_w3064_v = ~(v_w558_v & v_w851_v);
	assign v_w3905_v = ~(v_w3903_v & v_w3904_v);
	assign v_w4085_v = ~(v_w4084_v & v_w691_v);
	assign v_w6651_v = ~(v_w6649_v | v_w6650_v);
	assign v_w559_v = ~(v_s395_v & v_s473_v);
	assign v_w6762_v = ~(v_w1788_v & v_w895_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s218_v<=0;
	end
	else
	begin
	v_s218_v<=v_w231_v;
	end
	end
	assign v_w6303_v = ~(v_s207_v & v_w6278_v);
	assign v_w3441_v = ~(v_s361_v & v_w693_v);
	assign v_w2407_v = ~(v_w2406_v & v_w2327_v);
	assign v_w4209_v = ~(v_w4199_v & v_w4202_v);
	assign v_w5189_v = ~(v_w866_v | v_w1_v);
	assign v_w4131_v = ~(v_w692_v & v_w4130_v);
	assign v_w4121_v = v_w4117_v ^ v_w4120_v;
	assign v_w3919_v = ~(v_w3918_v & v_w3801_v);
	assign v_w1115_v = ~(v_w1329_v & v_w809_v);
	assign v_w7168_v = ~(v_w1386_v | v_w7117_v);
	assign v_w5202_v = ~(v_w5200_v | v_w5201_v);
	assign v_w3857_v = ~(v_w3735_v & v_w1131_v);
	assign v_w1667_v = ~(v_s335_v ^ v_w1666_v);
	assign v_w4123_v = ~(v_w887_v & v_w4116_v);
	assign v_w949_v = ~(v_w945_v | v_w830_v);
	assign v_w7769_v = ~(v_w847_v | v_w1782_v);
	assign v_w3581_v = ~(v_w3580_v & v_w3568_v);
	assign v_w5058_v = ~(v_w5055_v & v_w5057_v);
	assign v_w6477_v = ~(v_w6475_v & v_w6476_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s321_v<=0;
	end
	else
	begin
	v_s321_v<=v_w347_v;
	end
	end
	assign v_w2956_v = ~(v_w2951_v | v_w2955_v);
	assign v_w7728_v = ~(v_w7726_v & v_w7727_v);
	assign v_w2132_v = ~(v_w2130_v & v_w2131_v);
	assign v_w7302_v = ~(v_w7297_v & v_w7300_v);
	assign v_w7448_v = ~(v_w1134_v | v_w680_v);
	assign v_w1995_v = ~(v_w686_v | v_w1378_v);
	assign v_w795_v = ~(v_w1239_v & v_w751_v);
	assign v_w1574_v = ~(v_s247_v & v_w731_v);
	assign v_w1292_v = ~(v_w666_v & v_s442_v);
	assign v_w7802_v = ~(v_w654_v & v_w7801_v);
	assign v_w1762_v = ~(v_w1761_v);
	assign v_w6165_v = ~(v_w6151_v | v_w6164_v);
	assign v_w3376_v = ~(v_w3374_v & v_w3375_v);
	assign v_w5336_v = ~(v_w5331_v & v_w5335_v);
	assign v_w1447_v = ~(v_w1446_v | v_w1180_v);
	assign v_w7715_v = ~(v_w1783_v & v_w919_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s133_v<=0;
	end
	else
	begin
	v_s133_v<=v_w142_v;
	end
	end
	assign v_w1313_v = ~(v_w769_v ^ v_w1042_v);
	assign v_w7257_v = ~(v_w7252_v & v_w7256_v);
	assign v_w5593_v = ~(v_w675_v & v_w5442_v);
	assign v_w5377_v = ~(v_w683_v & v_w5376_v);
	assign v_w6545_v = v_s98_v ^ v_w1772_v;
	assign v_w7371_v = ~(v_w7369_v | v_w7370_v);
	assign v_w1404_v = ~(v_w1403_v);
	assign v_w2918_v = ~(v_w2915_v | v_w2917_v);
	assign v_w647_v = ~(v_w831_v ^ v_w945_v);
	assign v_w3659_v = ~(v_w3647_v & v_w3658_v);
	assign v_w838_v = ~(v_w1608_v & v_w1611_v);
	assign v_w3375_v = ~(v_w851_v & v_w2639_v);
	assign v_w5325_v = ~(v_w5125_v | v_w5034_v);
	assign v_w7380_v = ~(v_w687_v | v_w834_v);
	assign v_w1350_v = ~(v_w1348_v & v_w1349_v);
	assign v_w2199_v = ~(v_w2198_v & v_w2191_v);
	assign v_w4883_v = ~(v_w2347_v & v_w2870_v);
	assign v_w2109_v = ~(v_w1963_v | v_w1984_v);
	assign v_w5500_v = ~(v_w756_v | v_w2602_v);
	assign v_w3143_v = ~(v_w3142_v | v_w2606_v);
	assign v_w4107_v = ~(v_w4099_v | v_w4106_v);
	assign v_w8137_v = v_w8136_v ^ v_keyinput_50_v;
	assign v_w3611_v = ~(v_w3118_v);
	assign v_w5954_v = ~(v_w2053_v & v_w635_v);
	assign v_w6004_v = ~(v_w627_v & v_w2059_v);
	assign v_w6421_v = ~(v_w1440_v & v_w6019_v);
	assign v_w6554_v = ~(v_w6523_v & v_w6522_v);
	assign v_w776_v = ~(v_w710_v & v_s267_v);
	assign v_w3993_v = v_w3987_v & v_w3990_v;
	assign v_w7893_v = ~(v_s92_v & v_w7876_v);
	assign v_w3599_v = v_w3594_v & v_w3598_v;
	assign v_w4005_v = ~(v_w4003_v | v_w4004_v);
	assign v_w4423_v = ~(v_w3480_v | v_w4422_v);
	assign v_w2713_v = ~(v_w2709_v | v_w2712_v);
	assign v_w2663_v = ~(v_w2661_v & v_w2662_v);
	assign v_w8231_v = ~(v_w2326_v & v_w1131_v);
	assign v_w5006_v = ~(v_w674_v | v_w5005_v);
	assign v_w1341_v = ~(v_s78_v & v_w562_v);
	assign v_w7567_v = ~(v_w7564_v & v_w7566_v);
	assign v_w5770_v = ~(v_w1856_v | v_w2138_v);
	assign v_w4326_v = ~(v_w2784_v);
	assign v_w5822_v = ~(v_w2088_v ^ v_w2089_v);
	assign v_w1420_v = ~(v_s112_v & v_w562_v);
	assign v_w5977_v = ~(v_s303_v & v_w528_v);
	assign v_w5551_v = ~(v_w5037_v & v_w4424_v);
	assign v_w3102_v = ~(v_w3099_v & v_w3101_v);
	assign v_w7476_v = ~(v_w7348_v & v_w7475_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s459_v<=0;
	end
	else
	begin
	v_s459_v<=v_w512_v;
	end
	end
	assign v_w3693_v = ~(v_w3533_v);
	assign v_w1782_v = ~(v_w882_v & v_w1781_v);
	assign v_w747_v = ~(v_w1045_v & v_w996_v);
	assign v_w3986_v = ~(v_w755_v & v_w881_v);
	assign v_w6209_v = ~(v_s226_v & v_w1503_v);
	assign v_w2153_v = ~(v_s125_v | v_s171_v);
	assign v_w2142_v = ~(v_w2140_v & v_w2141_v);
	assign v_w1659_v = ~(v_w1654_v & v_w1658_v);
	assign v_w8216_v = v_w8215_v ^ v_keyinput_105_v;
	assign v_w120_v = ~(v_s486_v);
	assign v_w5124_v = ~(v_w5123_v);
	assign v_w7897_v = ~(v_s413_v & v_w7876_v);
	assign v_w525_v = ~(v_w6536_v & v_w6538_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s20_v<=0;
	end
	else
	begin
	v_s20_v<=v_w22_v;
	end
	end
	assign v_w5496_v = ~(v_w4662_v & v_w5495_v);
	assign v_w901_v = ~(v_w1453_v);
	assign v_w4373_v = ~(v_w4356_v | v_w4357_v);
	assign v_w5637_v = ~(v_w420_v & v_w2618_v);
	assign v_w5133_v = ~(v_w5132_v & v_w2257_v);
	assign v_w6190_v = ~(v_w6188_v & v_w6189_v);
	assign v_w2536_v = ~(v_w2534_v | v_w2535_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s384_v<=0;
	end
	else
	begin
	v_s384_v<=v_w430_v;
	end
	end
	assign v_w7640_v = ~(v_w7238_v | v_w7639_v);
	assign v_w6181_v = ~(v_w1514_v & v_w6154_v);
	assign v_w4853_v = ~(v_w4851_v | v_w4852_v);
	assign v_w5345_v = ~(v_w5342_v & v_w5344_v);
	assign v_w6093_v = ~(v_w6029_v | v_w6092_v);
	assign v_w6232_v = ~(v_w6230_v | v_w6231_v);
	assign v_w1877_v = ~(v_w1021_v & v_w1416_v);
	assign v_w4251_v = ~(v_s331_v ^ v_w2896_v);
	assign v_w6288_v = ~(v_s322_v & v_w6263_v);
	assign v_w4961_v = ~(v_w4959_v & v_w4960_v);
	assign v_w7504_v = ~(v_w7502_v | v_w7503_v);
	assign v_w7318_v = ~(v_w7313_v & v_w7316_v);
	assign v_w1750_v = ~(v_w1748_v & v_w1749_v);
	assign v_w5192_v = ~(v_w1703_v | v_w5145_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s254_v<=0;
	end
	else
	begin
	v_s254_v<=v_w269_v;
	end
	end
	assign v_w5279_v = ~(v_w3476_v | v_w4430_v);
	assign v_w3294_v = ~(v_w3290_v | v_w3293_v);
	assign v_w2990_v = ~(v_w2972_v | v_w2989_v);
	assign v_w7910_v = ~(v_w651_v & v_w7839_v);
	assign v_w6782_v = ~(v_s400_v & v_w656_v);
	assign v_w7914_v = ~(v_w651_v & v_w7849_v);
	assign v_w1797_v = ~(v_w660_v & v_w679_v);
	assign v_w906_v = ~(v_w3114_v & v_w2634_v);
	assign v_w897_v = ~(v_w2330_v);
	assign v_w172_v = ~(v_w5144_v & v_w5147_v);
	assign v_w2739_v = ~(v_w558_v & v_w2738_v);
	assign v_w6947_v = v_w953_v ^ v_w6909_v;
	assign v_w2330_v = v_w2329_v ^ v_s173_v;
	assign v_w2861_v = ~(v_w2856_v);
	assign v_w2987_v = ~(v_w1083_v | v_w617_v);
	assign v_w4299_v = ~(v_w4296_v & v_w4298_v);
	assign v_w2768_v = ~(v_s371_v & v_w2358_v);
	assign v_w1026_v = ~(v_w1127_v & v_w1128_v);
	assign v_w6856_v = ~(v_w1788_v & v_w1678_v);
	assign v_w987_v = ~(v_w1501_v & v_w1505_v);
	assign v_w6178_v = ~(v_w6176_v | v_w6177_v);
	assign v_w721_v = ~(v_w715_v & v_w345_v);
	assign v_w7247_v = ~(v_w1761_v & v_w680_v);
	assign v_w2736_v = ~(v_w2733_v | v_w2735_v);
	assign v_w7563_v = ~(v_w7560_v | v_w7562_v);
	assign v_w7367_v = ~(v_w1101_v | v_w680_v);
	assign v_w1265_v = ~(v_w1263_v & v_w1264_v);
	assign v_w249_v = ~(v_w7860_v & v_w7861_v);
	assign v_w1600_v = ~(v_w666_v & v_s206_v);
	assign v_w5292_v = v_w2253_v | v_w5134_v;
	assign v_w1584_v = ~(v_w1575_v & v_w1583_v);
	assign v_w1980_v = ~(v_w1979_v);
	assign v_w860_v = ~(v_w564_v & v_s32_v);
	assign v_w4645_v = v_w4417_v ^ v_w756_v;
	assign v_w5208_v = ~(v_w693_v | v_w2960_v);
	assign v_w1783_v = ~(v_w1782_v);
	assign v_w827_v = ~(v_w828_v | v_s283_v);
	assign v_w8205_v = v_w8204_v ^ v_keyinput_98_v;
	assign v_w3852_v = v_w3848_v | v_w3851_v;
	assign v_w7106_v = ~(v_w656_v & v_s35_v);
	assign v_w5592_v = ~(v_s105_v & v_w676_v);
	assign v_w7439_v = ~(v_w7372_v & v_w7438_v);
	assign v_w1172_v = v_s448_v ^ v_w1171_v;
	assign v_w3473_v = ~(v_s191_v & v_w699_v);
	assign v_w339_v = ~(v_w4988_v & v_w4993_v);
	assign v_w5918_v = ~(v_w2117_v & v_w997_v);
	assign v_w49_v = ~(v_w5604_v & v_w5605_v);
	assign v_w5543_v = ~(v_w3482_v | v_w2602_v);
	assign v_w3450_v = ~(v_w2358_v & v_s425_v);
	assign v_w4329_v = ~(v_s372_v & v_w4056_v);
	assign v_w726_v = ~(v_w724_v | v_w725_v);
	assign v_w7990_v = v_s467_v & v_s363_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s179_v<=0;
	end
	else
	begin
	v_s179_v<=v_w192_v;
	end
	end
	assign v_w7001_v = ~(v_w6999_v & v_w7000_v);
	assign v_w6391_v = ~(v_w5922_v & v_w6390_v);
	assign v_w7010_v = ~(v_w7008_v & v_w7009_v);
	assign v_w3589_v = ~(v_w3369_v | v_w1124_v);
	assign v_w1891_v = ~(v_w1811_v & v_w1890_v);
	assign v_w231_v = ~(v_w5162_v & v_w5163_v);
	assign v_w4476_v = ~(v_w4474_v | v_w4475_v);
	assign v_w3759_v = ~(v_w3757_v & v_w3758_v);
	assign v_w4466_v = ~(v_w3649_v | v_w4465_v);
	assign v_w1121_v = ~(v_w2300_v & v_w1277_v);
	assign v_w3185_v = ~(v_w3084_v & v_w3105_v);
	assign v_w6243_v = ~(v_s224_v & v_w6212_v);
	assign v_w962_v = ~(v_w961_v);
	assign v_w3982_v = ~(v_w3756_v & v_w3759_v);
	assign v_w5010_v = ~(v_w5008_v & v_w5009_v);
	assign v_w1531_v = ~(v_w1529_v & v_w1530_v);
	assign v_w1499_v = ~(v_w666_v & v_s223_v);
	assign v_w4568_v = ~(v_w3577_v | v_w4567_v);
	assign v_w4119_v = ~(v_w4108_v & v_w4111_v);
	assign v_w3868_v = v_w8072_v ^ v_keyinput_8_v;
	assign v_w6796_v = ~(v_w6789_v | v_w6795_v);
	assign v_w922_v = ~(v_w1826_v | v_w1852_v);
	assign v_w752_v = ~(v_in21_v ^ v_w1242_v);
	assign v_w6515_v = v_w6510_v | v_w6513_v;
	assign v_w6127_v = ~(v_w6125_v & v_w6126_v);
	assign v_w999_v = v_w1178_v & v_w484_v;
	assign v_w6706_v = ~(v_w6693_v | v_w6705_v);
	assign v_w1046_v = ~(v_in15_v & v_w1223_v);
	assign v_w4437_v = ~(v_w3482_v | v_w2264_v);
	assign v_w5984_v = v_w641_v ^ v_w642_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s151_v<=0;
	end
	else
	begin
	v_s151_v<=v_w160_v;
	end
	end
	assign v_w3785_v = ~(v_w3735_v | v_w2993_v);
	assign v_w119_v = ~(v_w5198_v & v_w5199_v);
	assign v_w1935_v = v_s68_v | v_s67_v;
	assign v_w7716_v = ~(v_w7714_v & v_w7715_v);
	assign v_w368_v = ~(v_w5953_v & v_w5956_v);
	assign v_w6555_v = ~(v_w6553_v & v_w6554_v);
	assign v_w1027_v = ~(v_w834_v);
	assign v_w7693_v = ~(v_w7660_v);
	assign v_w6665_v = ~(v_w6664_v & v_w6626_v);
	assign v_w6692_v = v_w6571_v | v_w1330_v;
	assign v_w87_v = ~(v_w7149_v & v_w7150_v);
	assign v_w3947_v = ~(v_w3944_v | v_w3946_v);
	assign v_w6602_v = ~(v_w1915_v);
	assign v_w5819_v = ~(v_w5817_v & v_w5818_v);
	assign v_w5542_v = ~(v_s191_v & v_w5386_v);
	assign v_w4619_v = ~(v_w4617_v | v_w4618_v);
	assign v_w7278_v = ~(v_w7276_v & v_w7277_v);
	assign v_w4806_v = ~(v_w4805_v | v_w4589_v);
	assign v_w7008_v = ~(v_s304_v & v_w656_v);
	assign v_w3507_v = ~(v_w2585_v & v_w2590_v);
	assign v_w2197_v = ~(v_s40_v & v_w2196_v);
	assign v_w2170_v = ~(v_s168_v | v_s165_v);
	assign v_w4362_v = v_w3017_v ^ v_s105_v;
	assign v_w8099_v = v_w8098_v ^ v_keyinput_25_v;
	assign v_w4174_v = ~(v_s229_v & v_w4153_v);
	assign v_w3411_v = ~(v_w3005_v & v_w2634_v);
	assign v_w1723_v = ~(v_w1719_v | v_w1722_v);
	assign v_w2994_v = ~(v_w2484_v & v_w2993_v);
	assign v_w7895_v = ~(v_s81_v & v_w7876_v);
	assign v_w6176_v = ~(v_w6029_v | v_w6175_v);
	assign v_w2613_v = ~(v_w2580_v & v_s293_v);
	assign v_w704_v = ~(v_w702_v & v_w703_v);
	assign v_w4849_v = ~(v_w4848_v | v_w4589_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s327_v<=0;
	end
	else
	begin
	v_s327_v<=v_w353_v;
	end
	end
	assign v_w498_v = ~(v_w6623_v & v_w6633_v);
	assign v_w5680_v = ~(v_s16_v & v_w695_v);
	assign v_w3100_v = ~(v_w3095_v);
	assign v_w1650_v = ~(v_w1648_v & v_w1649_v);
	assign v_w7796_v = ~(v_w654_v & v_w7795_v);
	assign v_w6126_v = ~(v_s273_v & v_w6099_v);
	assign v_w1805_v = ~(v_w1287_v | v_w1003_v);
	assign v_w3973_v = v_w8182_v ^ v_keyinput_84_v;
	assign v_w5337_v = ~(v_w683_v & v_w5336_v);
	assign v_w4044_v = v_s172_v & v_s256_v;
	assign v_w5886_v = ~(v_w1532_v | v_w2135_v);
	assign v_w447_v = ~(v_w7165_v & v_w7166_v);
	assign v_w2310_v = ~(v_w2294_v | v_w1542_v);
	assign v_w6035_v = ~(v_w6028_v | v_w6034_v);
	assign v_w7710_v = ~(v_w6987_v & v_w7709_v);
	assign v_w5313_v = ~(v_w683_v & v_w5312_v);
	assign v_w3027_v = ~(v_w3024_v & v_w3026_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s196_v<=0;
	end
	else
	begin
	v_s196_v<=v_w209_v;
	end
	end
	assign v_w5185_v = v_w5141_v & v_s93_v;
	assign v_w875_v = v_w874_v;
	assign v_w4688_v = ~(v_w4681_v & v_w4687_v);
	assign v_w3718_v = ~(v_w3594_v & v_w3717_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s130_v<=0;
	end
	else
	begin
	v_s130_v<=v_w139_v;
	end
	end
	assign v_w4810_v = v_s389_v & v_w674_v;
	assign v_w106_v = ~(v_w7891_v & v_w7892_v);
	assign v_w146_v = v_s137_v & v_w5134_v;
	assign v_w2527_v = ~(v_w2391_v | v_w538_v);
	assign v_w6139_v = ~(v_w1539_v | v_w6116_v);
	assign v_w6607_v = ~(v_w758_v & v_w6600_v);
	assign v_w7401_v = ~(v_w7399_v | v_w7400_v);
	assign v_w7629_v = ~(v_w912_v | v_w7628_v);
	assign v_w6273_v = v_w6268_v ^ v_w6272_v;
	assign v_w1358_v = ~(v_w1052_v & v_s81_v);
	assign v_w1166_v = ~(v_w1165_v & v_w461_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s189_v<=0;
	end
	else
	begin
	v_s189_v<=v_w202_v;
	end
	end
	assign v_w1949_v = ~(v_s48_v | v_s45_v);
	assign v_w6853_v = ~(v_w6851_v | v_w6852_v);
	assign v_w2650_v = ~(v_w2649_v & v_s379_v);
	assign v_w2686_v = ~(v_s385_v ^ v_w2657_v);
	assign v_w1285_v = ~(v_w1283_v & v_w1284_v);
	assign v_w364_v = ~(v_w7185_v & v_w7186_v);
	assign v_w2372_v = ~(v_w699_v & v_s230_v);
	assign v_w1146_v = ~(v_w6591_v & v_w6593_v);
	assign v_w5859_v = v_w5857_v ^ v_w5858_v;
	assign v_w3811_v = ~(v_w3809_v | v_w3810_v);
	assign v_w1872_v = ~(v_w1819_v & v_w1871_v);
	assign v_w6713_v = v_w1733_v ^ v_w1736_v;
	assign v_w1814_v = ~(v_w1813_v | v_w1384_v);
	assign v_w7847_v = ~(v_s419_v & v_w7742_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s407_v<=0;
	end
	else
	begin
	v_s407_v<=v_w456_v;
	end
	end
	assign v_w93_v = ~(v_w7153_v & v_w7154_v);
	assign v_w2533_v = ~(v_w2529_v ^ v_w2532_v);
	assign v_w6186_v = ~(v_w6185_v & v_w6020_v);
	assign v_w4759_v = ~(v_w1078_v | v_w2264_v);
	assign v_w2837_v = ~(v_w1099_v | v_w2836_v);
	assign v_w2618_v = ~(v_w2616_v & v_w2617_v);
	assign v_w5384_v = ~(v_w5381_v & v_w5383_v);
	assign v_w4987_v = ~(v_w4975_v & v_w4986_v);
	assign v_w6516_v = ~(v_w6514_v & v_w6515_v);
	assign v_w5761_v = ~(v_w5759_v & v_w5760_v);
	assign v_w5095_v = ~(v_w4527_v & v_w5085_v);
	assign v_w6664_v = v_w1899_v ^ v_w6659_v;
	assign v_w5614_v = ~(v_s19_v & v_w676_v);
	assign v_w2028_v = ~(v_w945_v | v_w2027_v);
	assign v_w6866_v = ~(v_w8222_v);
	assign v_w4659_v = ~(v_w4657_v & v_w4658_v);
	assign v_w7426_v = ~(v_w7411_v & v_w7425_v);
	assign v_w7242_v = ~(v_w687_v & v_w1762_v);
	assign v_w1180_v = ~(v_w870_v);
	assign v_w1190_v = v_s25_v ^ v_w1189_v;
	assign v_w5627_v = ~(v_w420_v & v_w2399_v);
	assign v_w6224_v = ~(v_w657_v & v_s306_v);
	assign v_w1050_v = ~(v_w1049_v & v_w1048_v);
	assign v_w7109_v = ~(v_s17_v | v_w7108_v);
	assign v_w887_v = ~(v_w885_v | v_w886_v);
	assign v_w1321_v = ~(v_w1317_v | v_w1320_v);
	assign v_w4219_v = ~(v_w4212_v & v_w4218_v);
	assign v_w2214_v = ~(v_s137_v | v_s136_v);
	assign v_w6590_v = ~(v_s453_v & v_w656_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s346_v<=0;
	end
	else
	begin
	v_s346_v<=v_w381_v;
	end
	end
	assign v_w8026_v = ~(v_w8024_v | v_w8025_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s216_v<=0;
	end
	else
	begin
	v_s216_v<=v_w229_v;
	end
	end
	assign v_w2207_v = ~(v_w2203_v | v_w2206_v);
	assign v_w1044_v = ~(v_w1043_v | v_w748_v);
	assign v_w7485_v = ~(v_w680_v & v_w1416_v);
	assign v_w426_v = ~(v_w3181_v & v_w3184_v);
	assign v_w6240_v = ~(v_w6239_v & v_w6020_v);
	assign v_w377_v = ~(v_s506_v);
	assign v_w41_v = ~(v_w7105_v & v_w7106_v);
	assign v_w865_v = ~(v_s171_v ^ v_w2231_v);
	assign v_w5033_v = ~(v_w5030_v | v_w5032_v);
	assign v_w6023_v = ~(v_w6019_v | v_w6022_v);
	assign v_w589_v = ~(v_in22_v | v_w1245_v);
	assign v_w6765_v = ~(v_w1710_v);
	assign v_w7930_v = ~(v_w527_v & v_w1100_v);
	assign v_w5156_v = ~(v_w1288_v | v_w5145_v);
	assign v_w3339_v = ~(v_w2607_v & v_w3338_v);
	assign v_w190_v = ~(v_w5410_v & v_w5417_v);
	assign v_w4018_v = ~(v_w3624_v | v_w4017_v);
	assign v_w8104_v = v_w8103_v ^ v_keyinput_28_v;
	assign v_w4518_v = ~(v_w4447_v | v_w4517_v);
	assign v_w1448_v = ~(v_w1052_v & v_s160_v);
	assign v_w3859_v = ~(v_w3857_v & v_w3858_v);
	assign v_w3482_v = ~(v_w3480_v);
	assign v_w2453_v = ~(v_w2349_v | v_w2452_v);
	assign v_w3114_v = v_w437_v ^ v_w3113_v;
	assign v_w1977_v = ~(v_s433_v | v_w1933_v);
	assign v_w2863_v = v_w2847_v ^ v_keyinput_53_v;
	assign v_w4229_v = ~(v_w4227_v & v_w4228_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s213_v<=0;
	end
	else
	begin
	v_s213_v<=v_w226_v;
	end
	end
	assign v_w4587_v = ~(v_w4585_v & v_w4586_v);
	assign v_w1211_v = ~(v_s82_v & v_w1192_v);
	assign v_w7638_v = ~(v_w7636_v & v_w7637_v);
	assign v_w337_v = ~(v_s499_v);
	assign v_w7600_v = ~(v_w1471_v | v_w7599_v);
	assign v_w7231_v = ~(v_w1579_v | v_w528_v);
	assign v_w5722_v = ~(v_w5720_v | v_w5721_v);
	assign v_w2673_v = ~(v_w8145_v);
	assign v_w2190_v = ~(v_s218_v & v_w531_v);
	assign v_w1571_v = ~(v_w665_v & v_s358_v);
	assign v_w8043_v = ~(v_w7987_v | v_w8042_v);
	assign v_w2081_v = v_w1999_v ^ v_w917_v;
	assign v_w4710_v = ~(v_w4708_v | v_w4709_v);
	assign v_w6345_v = ~(v_w6343_v ^ v_w6344_v);
	assign v_w597_v = ~(v_w2007_v | v_w1401_v);
	assign v_w1322_v = ~(v_w666_v & v_s416_v);
	assign v_w4233_v = ~(v_w4230_v | v_w4232_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s302_v<=0;
	end
	else
	begin
	v_s302_v<=v_w325_v;
	end
	end
	assign v_w2965_v = ~(v_w1088_v);
	assign v_w4382_v = ~(v_w3018_v | v_s105_v);
	assign v_w8193_v = v_w2603_v & v_w2622_v;
	assign v_w357_v = ~(v_w4943_v & v_w4956_v);
	assign v_w3862_v = ~(v_w3860_v & v_w3861_v);
	assign v_w489_v = ~(v_w6677_v & v_w6690_v);
	assign v_w5740_v = ~(v_w5738_v & v_w5739_v);
	assign v_w4183_v = ~(v_w4154_v & v_w4157_v);
	assign v_w8250_v = v_w8249_v ^ v_keyinput_125_v;
	assign v_w248_v = ~(v_w7691_v & v_w7692_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s397_v<=0;
	end
	else
	begin
	v_s397_v<=v_w446_v;
	end
	end
	assign v_w6081_v = ~(v_w6077_v ^ v_w6080_v);
	assign v_w914_v = ~(v_w3191_v & v_w1139_v);
	assign v_w3515_v = ~(v_w2585_v | v_w2590_v);
	assign v_w2644_v = ~(v_w2643_v & v_s328_v);
	assign v_w1618_v = ~(v_w870_v & v_w1617_v);
	assign v_w112_v = ~(v_w5594_v & v_w5595_v);
	assign v_w6977_v = ~(v_s308_v & v_w656_v);
	assign v_w3374_v = v_w8173_v ^ v_keyinput_77_v;
	assign v_w6637_v = ~(v_w884_v);
	assign v_w7550_v = ~(v_w7241_v | v_w7549_v);
	assign v_w5978_v = ~(v_w2137_v & v_w1100_v);
	assign v_w1621_v = ~(v_w874_v & v_s324_v);
	assign v_w4167_v = ~(v_w2554_v | v_w4041_v);
	assign v_w5355_v = ~(v_w2601_v & v_w2803_v);
	assign v_w2838_v = ~(v_w2830_v | v_w2835_v);
	assign v_w6634_v = ~(v_s441_v & v_w656_v);
	assign v_w5951_v = ~(v_w892_v & v_w1650_v);
	assign v_w4721_v = ~(v_w4717_v | v_w4720_v);
	assign v_w3486_v = ~(v_w565_v & v_s11_v);
	assign v_w581_v = ~(v_w579_v & v_w580_v);
	assign v_w1947_v = ~(v_w1943_v | v_w1946_v);
	assign v_w7507_v = ~(v_w679_v | v_w1337_v);
	assign v_w338_v = ~(v_w3328_v & v_w3330_v);
	assign v_w2459_v = ~(v_w2401_v | v_w2434_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s47_v<=0;
	end
	else
	begin
	v_s47_v<=v_w55_v;
	end
	end
	assign v_w1055_v = ~(v_w1106_v & v_w1107_v);
	assign v_w1834_v = ~(v_w8119_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s518_v<=0;
	end
	else
	begin
	v_s518_v<=v_w496_v;
	end
	end
	assign v_w5231_v = ~(v_s208_v & v_w5141_v);
	assign v_w3068_v = ~(v_w3063_v | v_w3067_v);
	assign v_w2221_v = ~(v_s129_v | v_s126_v);
	assign v_w2286_v = ~(v_w2151_v);
	assign v_w7976_v = ~(v_w527_v & v_w7253_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s4_v<=0;
	end
	else
	begin
	v_s4_v<=v_w4_v;
	end
	end
	assign v_w6182_v = ~(v_s288_v & v_w6155_v);
	assign v_w2258_v = ~(v_w2257_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s156_v<=0;
	end
	else
	begin
	v_s156_v<=v_w165_v;
	end
	end
	assign v_w3544_v = ~(v_w3540_v & v_w3543_v);
	assign v_w5344_v = ~(v_w5025_v | v_w5343_v);
	assign v_w3931_v = ~(v_w1079_v | v_w881_v);
	assign v_w4190_v = ~(v_w2799_v);
	assign v_w3964_v = v_w8124_v ^ v_keyinput_43_v;
	assign v_w2598_v = ~(v_w2597_v);
	assign v_w4285_v = ~(v_w2883_v ^ v_s119_v);
	assign v_w4163_v = ~(v_w4161_v & v_w4162_v);
	assign v_w5243_v = ~(v_s227_v & v_w5140_v);
	assign v_w3438_v = ~(v_w2956_v | v_w2606_v);
	assign v_w4050_v = ~(v_w4048_v & v_w4049_v);
	assign v_w2353_v = ~(v_w266_v | v_w531_v);
	assign v_w2901_v = ~(v_w2899_v & v_w2900_v);
	assign v_w6466_v = ~(v_w6437_v & v_w6465_v);
	assign v_w1186_v = ~(v_w666_v & v_s450_v);
	assign v_w6301_v = ~(v_w6029_v | v_w6300_v);
	assign v_w5506_v = ~(v_w4652_v & v_w5505_v);
	assign v_w3425_v = ~(v_s386_v & v_w693_v);
	assign v_w4332_v = ~(v_s369_v & v_w4315_v);
	assign v_w8080_v = v_w8079_v ^ v_keyinput_13_v;
	assign v_w1065_v = ~(v_w1064_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s292_v<=0;
	end
	else
	begin
	v_s292_v<=v_w312_v;
	end
	end
	assign v_w2440_v = ~(v_w2308_v | v_w2439_v);
	assign v_w3750_v = ~(v_w3745_v & v_w3748_v);
	assign v_w2021_v = ~(v_w608_v | v_w2020_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s413_v<=0;
	end
	else
	begin
	v_s413_v<=v_w464_v;
	end
	end
	assign v_w5263_v = ~(v_s87_v & v_w5141_v);
	assign v_w5171_v = ~(v_w5146_v & v_w1313_v);
	assign v_w4913_v = ~(v_w4911_v | v_w4912_v);
	assign v_w3194_v = ~(v_s430_v & v_w2358_v);
	assign v_w7540_v = ~(v_w7538_v & v_w7539_v);
	assign v_w6231_v = ~(v_w6018_v | v_w1490_v);
	assign v_w6550_v = ~(v_w6514_v & v_w6549_v);
	assign v_w1284_v = ~(v_w666_v & v_s446_v);
	assign v_w7353_v = ~(v_w680_v | v_w1095_v);
	assign v_w8037_v = ~(v_w7993_v | v_w8036_v);
	assign v_w7861_v = ~(v_w651_v & v_w7690_v);
	assign v_w5687_v = ~(v_w2137_v & v_w1135_v);
	assign v_w1796_v = ~(v_w1793_v | v_w1795_v);
	assign v_w1787_v = ~(v_w680_v | v_w660_v);
	assign v_w7202_v = ~(v_s318_v & v_w7112_v);
	assign v_w5829_v = ~(v_w662_v & v_w1435_v);
	assign v_w4350_v = ~(v_w4349_v & v_w692_v);
	assign v_w5350_v = ~(v_w5348_v & v_w5349_v);
	assign v_w2301_v = ~(v_w2300_v & v_w1524_v);
	assign v_w176_v = ~(v_s487_v);
	assign v_w2385_v = ~(v_w2384_v & v_w697_v);
	assign v_w7326_v = ~(v_w7321_v & v_w7324_v);
	assign v_w5605_v = ~(v_w5555_v & v_w5496_v);
	assign v_w767_v = ~(v_in10_v | v_w1207_v);
	assign v_w3963_v = ~(v_w3961_v | v_w3962_v);
	assign v_w7314_v = ~(v_w679_v | v_w1075_v);
	assign v_w4266_v = ~(v_w4244_v | v_w4243_v);
	assign v_w5781_v = ~(v_w5779_v & v_w5780_v);
	assign v_w8009_v = ~(v_s455_v | v_w8008_v);
	assign v_w7265_v = ~(v_w7261_v & v_w7264_v);
	assign v_w7103_v = ~(v_w7100_v | v_w7102_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s336_v<=0;
	end
	else
	begin
	v_s336_v<=v_w366_v;
	end
	end
	assign v_w1809_v = ~(v_w1311_v | v_w1065_v);
	assign v_w7719_v = ~(v_w6947_v | v_w1919_v);
	assign v_w7324_v = ~(v_w7322_v | v_w7323_v);
	assign v_w3085_v = ~(v_w1288_v | v_w2294_v);
	assign v_w1383_v = ~(v_s396_v & v_w562_v);
	assign v_w2103_v = ~(v_w723_v ^ v_w2102_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s183_v<=0;
	end
	else
	begin
	v_s183_v<=v_w196_v;
	end
	end
	assign v_w7944_v = ~(v_w527_v & v_w1453_v);
	assign v_w5137_v = ~(v_w531_v | v_w693_v);
	assign v_w1596_v = ~(v_w1512_v | v_w1595_v);
	assign v_w7486_v = ~(v_w679_v & v_w1021_v);
	assign v_w771_v = ~(v_in10_v ^ v_w1207_v);
	assign v_w4714_v = ~(v_w4711_v | v_w4713_v);
	assign v_w4327_v = ~(v_w4326_v | v_w4041_v);
	assign v_w1323_v = ~(v_w1321_v & v_w1322_v);
	assign v_w660_v = ~(v_w1374_v & v_w1786_v);
	assign v_w5333_v = ~(v_w2475_v & v_w5126_v);
	assign v_w668_v = ~(v_w667_v);
	assign v_w821_v = ~(v_w564_v & v_s93_v);
	assign v_w6776_v = ~(v_w8143_v);
	assign v_w2836_v = ~(v_w2830_v ^ v_w2835_v);
	assign v_w1899_v = ~(v_w1810_v | v_w1898_v);
	assign v_w6161_v = v_w1514_v ^ v_w6160_v;
	assign v_w1173_v = v_s375_v | v_s374_v;
	assign v_w2007_v = ~(v_w723_v ^ v_w847_v);
	assign v_w7235_v = ~(v_s477_v & v_s475_v);
	assign v_w1656_v = ~(v_w1650_v);
	assign v_w3072_v = ~(v_w3070_v & v_w3071_v);
	assign v_w2433_v = ~(v_w2409_v | v_w2432_v);
	assign v_w1687_v = ~(v_w1454_v & v_w1686_v);
	assign v_w3330_v = ~(v_w3329_v & v_w3126_v);
	assign v_w1806_v = ~(v_w1003_v);
	assign v_w7203_v = ~(v_w1474_v | v_w528_v);
	assign v_w1998_v = ~(v_w1997_v | v_w1309_v);
	assign v_w7089_v = ~(v_w7088_v & v_w6639_v);
	assign v_w6669_v = ~(v_w6667_v & v_w6668_v);
	assign v_w6254_v = ~(v_w6252_v & v_w6253_v);
	assign v_w4128_v = ~(v_w4101_v & v_w4103_v);
	assign v_w4585_v = ~(v_w4584_v & v_w878_v);
	assign v_w7270_v = ~(v_w1311_v & v_w680_v);
	assign v_w5166_v = ~(v_w5164_v | v_w5165_v);
	assign v_w2556_v = ~(v_w2549_v | v_w2555_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s513_v<=0;
	end
	else
	begin
	v_s513_v<=v_w424_v;
	end
	end
	assign v_w7571_v = ~(v_w7563_v & v_w7570_v);
	assign v_w4342_v = ~(v_w692_v & v_w4341_v);
	assign v_w4353_v = ~(v_w2756_v & v_w887_v);
	assign v_w6501_v = ~(v_w6500_v & v_w6020_v);
	assign v_w2851_v = ~(v_s326_v ^ v_w2850_v);
	assign v_w8035_v = ~(v_w7995_v | v_w8034_v);
	assign v_w1619_v = ~(v_w1052_v & v_s205_v);
	assign v_w5162_v = ~(v_w5160_v | v_w5161_v);
	assign v_w6274_v = ~(v_w6029_v | v_w6273_v);
	assign v_w7967_v = ~(v_s22_v & v_w2143_v);
	assign v_w3684_v = v_w3683_v ^ v_w866_v;
	assign v_w6958_v = ~(v_w6956_v & v_w6957_v);
	assign v_w8042_v = ~(v_w7988_v | v_w8041_v);
	assign v_w8082_v = v_in27_v | v_w1262_v;
	assign v_w6169_v = ~(v_s234_v & v_w889_v);
	assign v_w1939_v = ~(v_w1935_v | v_w1938_v);
	assign v_w634_v = ~(v_w2051_v & v_w2053_v);
	assign v_w5045_v = ~(v_w2378_v | v_w2370_v);
	assign v_w4663_v = ~(v_w4655_v & v_w4662_v);
	assign v_w3108_v = ~(v_w1139_v & v_w3107_v);
	assign v_w5692_v = ~(v_w5688_v | v_w5691_v);
	assign v_w2780_v = ~(v_w2779_v & v_w384_v);
	assign v_w4002_v = ~(v_w3605_v & v_w881_v);
	assign v_w2955_v = ~(v_w2953_v & v_w2954_v);
	assign v_w7245_v = ~(v_w1769_v);
	assign v_w6215_v = ~(v_s304_v & v_w1503_v);
	assign v_w1401_v = ~(v_w1399_v & v_w1400_v);
	assign v_w7473_v = ~(v_w7357_v & v_w7472_v);
	assign v_w8105_v = ~(v_w1129_v & v_w1130_v);
	assign v_w1372_v = ~(v_w1370_v & v_w1371_v);
	assign v_w7992_v = v_s466_v & v_s353_v;
	assign v_w3219_v = ~(v_w3217_v & v_w3218_v);
	assign v_w5373_v = ~(v_w2601_v & v_w2861_v);
	assign v_w1365_v = ~(v_w1364_v);
	assign v_w537_v = ~(v_w539_v);
	assign v_o3_v = v_w8047_v ^ v_w8054_v;
	assign v_w148_v = v_s139_v & v_w5134_v;
	assign v_w7148_v = v_w7113_v & v_s78_v;
	assign v_w5921_v = ~(v_w5919_v | v_w5920_v);
	assign v_w6318_v = ~(v_s197_v ^ v_w6317_v);
	assign v_w2908_v = ~(v_w2905_v | v_w2907_v);
	assign v_w1975_v = ~(v_w1973_v | v_w1974_v);
	assign v_w4757_v = ~(v_w3031_v & v_w2347_v);
	assign v_w354_v = ~(v_w3158_v & v_w3159_v);
	assign v_w3535_v = ~(v_w2910_v & v_w2916_v);
	assign v_w7299_v = ~(v_w1726_v | v_w680_v);
	assign v_w7892_v = ~(v_w651_v & v_w7783_v);
	assign v_w3783_v = ~(v_w3781_v | v_w3782_v);
	assign v_w1849_v = ~(v_w1848_v & v_w790_v);
	assign v_w5123_v = ~(v_w2259_v & v_w879_v);
	assign v_w3427_v = ~(v_w2635_v | v_w2667_v);
	assign v_w573_v = ~(v_w1571_v & v_w1572_v);
	assign v_w6321_v = ~(v_w6299_v & v_w6295_v);
	assign v_w5460_v = ~(v_w5456_v & v_w5459_v);
	assign v_w4779_v = ~(v_w2448_v & v_w2761_v);
	assign v_w826_v = ~(v_w2054_v | v_w1126_v);
	assign v_w1607_v = v_w8146_v ^ v_keyinput_56_v;
	assign v_w4041_v = ~(v_w887_v);
	assign v_w873_v = v_w871_v | v_w872_v;
	assign v_w4686_v = ~(v_w4685_v | v_w4589_v);
	assign v_w329_v = ~(v_w6989_v & v_w6994_v);
	assign v_w2119_v = ~(v_w680_v & v_w1968_v);
	assign v_w2174_v = v_s275_v | v_s249_v;
	assign v_w3677_v = ~(v_w3627_v & v_w3676_v);
	assign v_w2642_v = ~(v_w2641_v & v_s313_v);
	assign v_w3772_v = ~(v_w3172_v & v_w881_v);
	assign v_w2587_v = ~(v_w2576_v & v_w2586_v);
	assign v_w1457_v = ~(v_w1455_v & v_w1456_v);
	assign v_w7328_v = ~(v_w679_v | v_w1436_v);
	assign v_w4336_v = ~(v_w4329_v & v_w4335_v);
	assign v_w7766_v = ~(v_w654_v & v_w7765_v);
	assign v_w2130_v = ~(v_w2125_v & v_w2129_v);
	assign v_w6292_v = v_w8110_v ^ v_keyinput_34_v;
	assign v_w8133_v = v_w8132_v ^ v_keyinput_48_v;
	assign v_w2114_v = ~(v_w2104_v & v_w2113_v);
	assign v_w2495_v = ~(v_w2493_v | v_w2494_v);
	assign v_w3315_v = ~(v_w2525_v ^ v_w2533_v);
	assign v_w706_v = v_w2155_v & v_w959_v;
	assign v_w1430_v = ~(v_w875_v & v_s354_v);
	assign v_w5454_v = ~(v_w4743_v & v_w5453_v);
	assign v_w3377_v = ~(v_w2635_v | v_w3056_v);
	assign v_w3807_v = ~(v_w3805_v | v_w3806_v);
	assign v_w5079_v = ~(v_w5077_v & v_w5078_v);
	assign v_w7085_v = ~(v_w1798_v & v_w602_v);
	assign v_w5861_v = ~(v_w2117_v & v_w1817_v);
	assign v_w5330_v = ~(v_w2296_v | v_w2602_v);
	assign v_w1361_v = ~(v_w875_v & v_s409_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s451_v<=0;
	end
	else
	begin
	v_s451_v<=v_w504_v;
	end
	end
	assign v_w2608_v = ~(v_w2607_v & v_w2367_v);
	assign v_w3882_v = ~(v_w3880_v | v_w3881_v);
	assign v_w75_v = v_s67_v & v_w7107_v;
	assign v_w3467_v = ~(v_w3465_v & v_w3466_v);
	assign v_w3268_v = ~(v_w3264_v | v_w3267_v);
	assign v_w7672_v = ~(v_w7087_v & v_w7671_v);
	assign v_w885_v = ~(v_s1_v & v_w694_v);
	assign v_w5952_v = ~(v_w5950_v & v_w5951_v);
	assign v_w107_v = ~(v_w7953_v & v_w7954_v);
	assign v_w5521_v = ~(v_w5520_v | v_w4611_v);
	assign v_w5088_v = ~(v_w5080_v & v_w5087_v);
	assign v_w5556_v = ~(v_s258_v & v_w676_v);
	assign v_w4897_v = ~(v_w4896_v & v_w673_v);
	assign v_w695_v = v_w693_v | v_w694_v;
	assign v_w5361_v = ~(v_w683_v & v_w5360_v);
	assign v_w5038_v = ~(v_w5036_v & v_w5037_v);
	assign v_w3880_v = ~(v_w2590_v | v_w3735_v);
	assign v_w724_v = ~(v_w1624_v | v_w1823_v);
	assign v_w1136_v = ~(v_w701_v ^ v_s164_v);
	assign v_w909_v = v_w365_v & v_w367_v;
	assign v_w4904_v = ~(v_w2342_v | v_w4903_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s145_v<=0;
	end
	else
	begin
	v_s145_v<=v_w154_v;
	end
	end
	assign v_w2974_v = ~(v_w2358_v & v_s369_v);
	assign v_w1602_v = v_s321_v ^ v_w1152_v;
	assign v_w6968_v = ~(v_w6964_v & v_w6967_v);
	assign v_w4214_v = ~(v_s212_v | v_w4190_v);
	assign v_w2749_v = v_s379_v ^ v_w2649_v;
	assign v_w6939_v = ~(v_w6592_v & v_w1632_v);
	assign v_w7192_v = ~(v_w1646_v | v_w7117_v);
	assign v_o12_v = ~(v_w8027_v ^ v_w8028_v);
	assign v_w5576_v = ~(v_s202_v & v_w676_v);
	assign v_w6472_v = v_s89_v ^ v_w6457_v;
	assign v_w7262_v = ~(v_w687_v | v_w1806_v);
	assign v_w3422_v = ~(v_w2547_v ^ v_w3421_v);
	assign v_w1458_v = ~(v_w666_v & v_s194_v);
	assign v_w2080_v = ~(v_w2077_v | v_w2079_v);
	assign v_w3902_v = ~(v_w3900_v & v_w3901_v);
	assign v_w1153_v = v_s321_v | v_w1152_v;
	assign v_w6576_v = ~(v_w6574_v & v_w6575_v);
	assign v_w3412_v = ~(v_s1_v | v_w314_v);
	assign v_w7511_v = ~(v_w7505_v | v_w7510_v);
	assign v_w7543_v = v_w7537_v & v_w7540_v;
	assign v_w749_v = ~(v_in21_v | v_w1242_v);
	assign v_w7298_v = ~(v_w679_v | v_w998_v);
	assign v_w5034_v = ~(v_w8068_v);
	assign v_w5367_v = ~(v_w5365_v | v_w5366_v);
	assign v_w4578_v = ~(v_w1008_v);
	assign v_w6386_v = ~(v_w6384_v & v_w6385_v);
	assign v_w1832_v = ~(v_w729_v & v_w596_v);
	assign v_w3514_v = ~(v_w3506_v & v_w3513_v);
	assign v_w8238_v = ~(v_w4458_v & v_w4469_v);
	assign v_w6026_v = ~(v_w664_v & v_s454_v);
	assign v_w5520_v = ~(v_w4604_v | v_w5123_v);
	assign v_w1090_v = ~(v_w1427_v | v_w808_v);
	assign v_w3092_v = ~(v_w2660_v & v_w697_v);
	assign v_w3707_v = ~(v_w3691_v | v_w3706_v);
	assign v_w3351_v = ~(v_w3349_v | v_w3350_v);
	assign v_w8050_v = ~(v_w7980_v & v_w8049_v);
	assign v_w4094_v = ~(v_w692_v & v_w4093_v);
	assign v_w6614_v = ~(v_w1172_v | v_w6571_v);
	assign v_w5256_v = ~(v_w1561_v | v_w5145_v);
	assign v_w5046_v = ~(v_w5044_v | v_w5045_v);
	assign v_w6068_v = ~(v_w664_v & v_s456_v);
	assign v_w673_v = ~(v_w2256_v & v_w2261_v);
	assign v_w2351_v = ~(v_w2350_v);
	assign v_w7081_v = ~(v_w1833_v | v_w1836_v);
	assign v_w1482_v = ~(v_w1480_v & v_w1481_v);
	assign v_w5823_v = ~(v_w2113_v & v_w5822_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s149_v<=0;
	end
	else
	begin
	v_s149_v<=v_w158_v;
	end
	end
	assign v_w6220_v = ~(v_w6219_v & v_w6020_v);
	assign v_w4818_v = ~(v_w967_v | v_w2264_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s334_v<=0;
	end
	else
	begin
	v_s334_v<=v_w362_v;
	end
	end
	assign v_w413_v = ~(v_w4324_v & v_w4325_v);
	assign v_w4632_v = ~(v_w4630_v | v_w4631_v);
	assign v_w3802_v = ~(v_w3732_v | v_w2937_v);
	assign v_w6203_v = ~(v_w6200_v ^ v_w6202_v);
	assign v_w1714_v = ~(v_w1385_v | v_w1713_v);
	assign v_w4789_v = ~(v_w864_v | v_w2264_v);
	assign v_w5528_v = ~(v_w5037_v & v_w4531_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s17_v<=0;
	end
	else
	begin
	v_s17_v<=v_w18_v;
	end
	end
	assign v_w682_v = ~(v_w2245_v | v_w2252_v);
	assign v_w3537_v = ~(v_w2926_v | v_w2935_v);
	assign v_w6506_v = ~(v_w6501_v & v_w6505_v);
	assign v_w5306_v = ~(v_w2326_v | v_w2602_v);
	assign v_w6786_v = ~(v_w6784_v | v_w6785_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s190_v<=0;
	end
	else
	begin
	v_s190_v<=v_w203_v;
	end
	end
	assign v_w114_v = ~(v_w5590_v & v_w5591_v);
	assign v_w98_v = ~(v_w7947_v & v_w7948_v);
	assign v_w5679_v = ~(v_w4082_v & v_w3485_v);
	assign v_w1756_v = ~(v_w1754_v & v_w1755_v);
	assign v_w407_v = ~(v_w4862_v & v_w4879_v);
	assign v_w7977_v = ~(v_s4_v & v_w2143_v);
	assign v_w4672_v = ~(v_w4670_v | v_w4671_v);
	assign v_w3795_v = ~(v_w2965_v & v_w3732_v);
	assign v_w2785_v = ~(v_w569_v & v_w2784_v);
	assign v_w7051_v = ~(v_w1788_v & v_w602_v);
	assign v_w6936_v = ~(v_w6935_v | v_w6640_v);
	assign v_w3200_v = ~(v_w3199_v | v_w2620_v);
	assign v_w3558_v = ~(v_w1079_v | v_w3012_v);
	assign v_w5626_v = ~(v_s242_v & v_w695_v);
	assign v_w1566_v = ~(v_s158_v & v_w870_v);
	assign v_w356_v = ~(v_w3383_v & v_w3391_v);
	assign v_w655_v = v_w1140_v | v_w1141_v;
	assign v_w6821_v = ~(v_w1816_v | v_w1797_v);
	assign v_w812_v = ~(v_w810_v | v_w811_v);
	assign v_w69_v = v_s61_v & v_w7107_v;
	assign v_w5037_v = ~(v_w4863_v);
	assign v_w2977_v = ~(v_w2976_v & v_w697_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s398_v<=0;
	end
	else
	begin
	v_s398_v<=v_w447_v;
	end
	end
	assign v_w187_v = ~(v_w5289_v | v_w5290_v);
	assign v_w2476_v = ~(v_w2458_v & v_w2475_v);
	assign v_w3209_v = ~(v_w3205_v | v_w3208_v);
	assign v_w6413_v = ~(v_w6029_v | v_w6412_v);
	assign v_w8064_v = v_w8063_v ^ v_keyinput_1_v;
	assign v_w510_v = ~(v_w6110_v & v_w6122_v);
	assign v_w861_v = ~(v_w2300_v & v_w1313_v);
	assign v_w849_v = ~(v_w1053_v | v_w1054_v);
	assign v_w3395_v = v_w2511_v ^ v_w2519_v;
	assign v_w7931_v = ~(v_s216_v & v_w6015_v);
	assign v_w4615_v = ~(v_w4600_v | v_w4614_v);
	assign v_w1308_v = ~(v_w666_v & v_s417_v);
	assign v_w7969_v = ~(v_s18_v & v_w2143_v);
	assign v_w5225_v = ~(v_w5145_v | v_w1628_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s442_v<=0;
	end
	else
	begin
	v_s442_v<=v_w494_v;
	end
	end
	assign v_w3172_v = ~(v_w2738_v);
	assign v_w1695_v = ~(v_w875_v & v_s400_v);
	assign v_w6013_v = ~(v_w5685_v | v_w663_v);
	assign v_w6370_v = ~(v_s344_v & v_w1465_v);
	assign v_w3371_v = ~(v_w3368_v | v_w3370_v);
	assign v_w609_v = v_w2015_v & v_w1830_v;
	assign v_w2743_v = ~(v_w2484_v & v_w2738_v);
	assign v_w7558_v = ~(v_w790_v | v_w979_v);
	assign v_w3661_v = ~(v_w3644_v & v_w3660_v);
	assign v_w1962_v = ~(v_s47_v | v_w1961_v);
	assign v_w3937_v = ~(v_w3777_v | v_w3929_v);
	assign v_w8032_v = ~(v_w8030_v | v_w8031_v);
	assign v_o6_v = v_w8041_v ^ v_w8057_v;
	assign v_w6465_v = ~(v_w6433_v & v_w6438_v);
	assign v_w6191_v = ~(v_w6187_v ^ v_w6190_v);
	assign v_w5957_v = ~(v_w2117_v & v_w2016_v);
	assign v_w2911_v = ~(v_w558_v & v_w2910_v);
	assign v_w3163_v = ~(v_w2317_v & v_w2639_v);
	assign v_w4561_v = ~(v_w3552_v & v_w4560_v);
	assign v_w5565_v = ~(v_w675_v & v_w5327_v);
	assign v_w839_v = ~(v_w837_v | v_w838_v);
	assign v_w2222_v = ~(v_w2220_v & v_w2221_v);
	assign v_w5301_v = ~(v_w5299_v & v_w5300_v);
	assign v_w3690_v = ~(v_w3570_v);
	assign v_w4553_v = ~(v_w3492_v | v_w4552_v);
	assign v_w3900_v = ~(v_w2916_v & v_w3732_v);
	assign v_w85_v = ~(v_w5600_v & v_w5601_v);
	assign v_w57_v = v_s49_v & v_w7107_v;
	assign v_w3006_v = ~(v_w3005_v & v_w697_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s348_v<=0;
	end
	else
	begin
	v_s348_v<=v_w383_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s419_v<=0;
	end
	else
	begin
	v_s419_v<=v_w470_v;
	end
	end
	assign v_w4257_v = v_w4054_v & v_s353_v;
	assign v_w5135_v = ~(v_w990_v | v_w2350_v);
	assign v_w7189_v = ~(v_w7187_v | v_w7188_v);
	assign v_w3403_v = ~(v_s1_v | v_w425_v);
	assign v_w1219_v = ~(v_w612_v & v_s396_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s60_v<=0;
	end
	else
	begin
	v_s60_v<=v_w68_v;
	end
	end
	assign v_w2032_v = ~(v_w723_v ^ v_w920_v);
	assign v_w2549_v = ~(v_w1506_v | v_w2294_v);
	assign v_w1389_v = ~(v_s374_v | v_w1388_v);
	assign v_w8153_v = v_w8152_v ^ v_keyinput_61_v;
	assign v_w1825_v = ~(v_w1824_v | v_w1632_v);
	assign v_w4637_v = ~(v_w4635_v & v_w4636_v);
	assign v_w2821_v = ~(v_s208_v & v_w565_v);
	assign v_w1581_v = ~(v_w613_v & v_w1580_v);
	assign v_w2685_v = ~(v_w2683_v & v_w2684_v);
	assign v_w6305_v = v_s205_v ^ v_w1626_v;
	assign v_w4419_v = ~(v_w871_v | v_w4418_v);
	assign v_w858_v = v_w912_v | v_w913_v;
	assign v_w2365_v = ~(v_w2360_v | v_w2364_v);
	assign v_w4832_v = ~(v_w2447_v & v_w2993_v);
	assign v_w3580_v = ~(v_w3578_v & v_w3579_v);
	assign v_w2355_v = v_w593_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s232_v<=0;
	end
	else
	begin
	v_s232_v<=v_w245_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s210_v<=0;
	end
	else
	begin
	v_s210_v<=v_w223_v;
	end
	end
	assign v_w566_v = ~(v_w1541_v | v_w1543_v);
	assign v_w854_v = ~(v_w856_v | v_w857_v);
	assign v_w1079_v = ~(v_w864_v);
	assign v_w6034_v = v_w8230_v ^ v_keyinput_114_v;
	assign v_w6327_v = v_w6322_v ^ v_w6326_v;
	assign v_w6142_v = ~(v_s236_v & v_w889_v);
	assign v_w5828_v = ~(v_s475_v | v_w377_v);
	assign v_w7791_v = ~(v_s91_v & v_w7742_v);
	assign v_w7276_v = ~(v_w687_v & v_w1323_v);
	assign v_w4760_v = ~(v_w4758_v | v_w4759_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s198_v<=0;
	end
	else
	begin
	v_s198_v<=v_w211_v;
	end
	end
	assign v_w92_v = ~(v_w5662_v & v_w5663_v);
	assign v_w3575_v = ~(v_w3077_v | v_w3574_v);
	assign v_w7463_v = v_w7459_v | v_w7462_v;
	assign v_w1655_v = ~(v_w1642_v);
	assign v_w2063_v = v_w2060_v | v_w1418_v;
	assign v_w7378_v = ~(v_w7376_v | v_w7377_v);
	assign v_w3836_v = ~(v_w3832_v & v_w3835_v);
	assign v_w6047_v = ~(v_w713_v | v_w396_v);
	assign v_w7670_v = ~(v_w7660_v & v_w7088_v);
	assign v_w1721_v = ~(v_w875_v & v_s405_v);
	assign v_w5335_v = ~(v_w2450_v | v_w5334_v);
	assign v_w2952_v = v_w401_v ^ v_w2646_v;
	assign v_w2416_v = ~(v_w2412_v | v_w2415_v);
	assign v_w4073_v = v_s266_v ^ v_w2321_v;
	assign v_w3597_v = ~(v_w3100_v | v_w3087_v);
	assign v_w269_v = ~(v_w5298_v & v_w5304_v);
	assign v_w4724_v = ~(v_w4722_v | v_w4723_v);
	assign v_w1390_v = ~(v_w1389_v | v_w8_v);
	assign v_w3634_v = v_w3556_v & v_w3563_v;
	assign v_w6025_v = ~(v_w6024_v & v_s477_v);
	assign v_w3773_v = ~(v_w3771_v & v_w3772_v);
	assign v_w905_v = ~(v_w903_v & v_w904_v);
	assign v_w1972_v = ~(v_w1971_v);
	assign v_w918_v = ~(v_w917_v);
	assign v_w3000_v = ~(v_w2998_v | v_w2999_v);
	assign v_w8033_v = ~(v_w7997_v | v_w8032_v);
	assign v_w6708_v = ~(v_w1787_v & v_w1362_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s120_v<=0;
	end
	else
	begin
	v_s120_v<=v_w129_v;
	end
	end
	assign v_w6247_v = ~(v_w6240_v & v_w6246_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s470_v<=0;
	end
	else
	begin
	v_s470_v<=v_w523_v;
	end
	end
	assign v_w2439_v = ~(v_w2391_v);
	assign v_w5056_v = ~(v_w2459_v ^ v_w2468_v);
	assign v_o20_v = v_s259_v ^ v_s454_v;
	assign v_w2574_v = ~(v_w565_v & v_s309_v);
	assign v_w7359_v = ~(v_w687_v | v_w1655_v);
	assign v_w7788_v = ~(v_w7786_v | v_w7787_v);
	assign v_w6373_v = v_w1667_v ^ v_w6372_v;
	assign v_w1272_v = v_in18_v ^ v_w1232_v;
	assign v_w572_v = ~(v_w570_v | v_w571_v);
	assign v_w518_v = ~(v_w6319_v & v_w6340_v);
	assign v_w355_v = ~(v_s501_v);
	assign v_w3924_v = ~(v_w3917_v | v_w3923_v);
	assign v_w3883_v = ~(v_w2575_v | v_w3731_v);
	assign v_w222_v = ~(v_w5362_v & v_w5369_v);
	assign v_w2256_v = ~(v_w682_v & v_w2255_v);
	assign v_w2012_v = ~(v_w723_v ^ v_w834_v);
	assign v_w2361_v = v_w696_v;
	assign v_w2260_v = ~(v_w8113_v);
	assign v_w5120_v = ~(v_w2265_v | v_w2343_v);
	assign v_w5158_v = ~(v_w5156_v | v_w5157_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s95_v<=0;
	end
	else
	begin
	v_s95_v<=v_w103_v;
	end
	end
	assign v_w4673_v = v_w753_v ^ v_w4416_v;
	assign v_w5752_v = ~(v_w5748_v | v_w5751_v);
	assign v_w4993_v = ~(v_w4991_v | v_w4992_v);
	assign v_w4301_v = ~(v_w2884_v & v_s119_v);
	assign v_w4265_v = ~(v_w2896_v | v_s200_v);
	assign v_w2082_v = ~(v_w2080_v | v_w2081_v);
	assign v_w3987_v = ~(v_w3985_v & v_w3986_v);
	assign v_w5503_v = ~(v_w5501_v & v_w5502_v);
	assign v_w2078_v = ~(v_w2075_v ^ v_w2076_v);
	assign v_w1752_v = ~(v_w1188_v & v_w893_v);
	assign v_w588_v = ~(v_w587_v | v_s300_v);
	assign v_w3850_v = ~(v_w2309_v & v_w3731_v);
	assign v_w3789_v = ~(v_w1083_v | v_w3735_v);
	assign v_w2631_v = ~(v_w2263_v & v_s1_v);
	assign v_w7091_v = ~(v_w7090_v & v_w655_v);
	assign v_w212_v = ~(v_w5378_v & v_w5385_v);
	assign v_w2726_v = ~(v_w558_v & v_w820_v);
	assign v_w4872_v = ~(v_w4870_v & v_w4871_v);
	assign v_w4652_v = ~(v_w4650_v | v_w4651_v);
	assign v_w3766_v = ~(v_w3764_v & v_w3765_v);
	assign v_w1717_v = ~(v_s95_v & v_w562_v);
	assign v_w6352_v = ~(v_w6350_v | v_w6351_v);
	assign v_w5360_v = v_w4979_v | v_w5359_v;
	assign v_w3423_v = ~(v_w3422_v & v_w3126_v);
	assign v_w6748_v = ~(v_w6747_v & v_w6626_v);
	assign v_w7315_v = ~(v_w1699_v | v_w680_v);
	assign v_w561_v = ~(v_w612_v | v_w613_v);
	assign v_w972_v = ~(v_w1022_v & v_w1023_v);
	assign v_w1368_v = ~(v_w870_v & v_w1367_v);
	assign v_w4621_v = ~(v_w8207_v);
	assign v_w3856_v = ~(v_w3854_v & v_w3855_v);
	assign v_w3778_v = ~(v_w3735_v | v_w2791_v);
	assign v_w6494_v = ~(v_w6490_v ^ v_w6493_v);
	assign v_w4893_v = ~(v_w4891_v & v_w4892_v);
	assign v_w1098_v = ~(v_w2807_v | v_w581_v);
	assign v_w2538_v = ~(v_w2296_v | v_w617_v);
	assign v_w1491_v = v_w1490_v | v_w1374_v;
	assign v_w1114_v = ~(v_w1112_v | v_w1113_v);
	assign v_w6150_v = ~(v_w664_v & v_s459_v);
	assign v_w1816_v = ~(v_w1401_v);
	assign v_w5872_v = ~(v_w892_v & v_w1066_v);
	assign v_w2487_v = ~(v_w2482_v | v_w2486_v);
	assign v_w331_v = ~(v_w6976_v & v_w6977_v);
	assign v_w2057_v = v_w1453_v ^ v_w900_v;
	assign v_w3060_v = ~(v_w3058_v & v_w3059_v);
	assign v_w5494_v = ~(v_w5123_v | v_w4660_v);
	assign v_w1413_v = ~(v_w1412_v | v_w1180_v);
	assign v_w3673_v = ~(v_w3631_v & v_w3672_v);
	assign v_w3010_v = ~(v_w2358_v & v_s391_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s392_v<=0;
	end
	else
	begin
	v_s392_v<=v_w441_v;
	end
	end
	assign v_w6430_v = ~(v_s114_v ^ v_w6429_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s521_v<=0;
	end
	else
	begin
	v_s521_v<=v_w532_v;
	end
	end
	assign v_w3266_v = ~(v_w3109_v & v_w2761_v);
	assign v_w2916_v = ~(v_w2901_v);
	assign v_w4231_v = ~(v_w4226_v & v_w4229_v);
	assign v_w3316_v = v_w8069_v ^ v_keyinput_4_v;
	assign v_w4514_v = ~(v_w8141_v);
	assign v_w312_v = ~(v_w3284_v & v_w3285_v);
	assign v_w3096_v = ~(v_w3095_v | v_w993_v);
	assign v_w7214_v = ~(v_s298_v & v_w7112_v);
	assign v_w5741_v = v_w2046_v ^ v_w2048_v;
	assign v_w177_v = ~(v_w5291_v & v_w5292_v);
	assign v_w5143_v = v_w544_v & v_s1_v;
	assign v_w964_v = ~(v_w963_v);
	assign v_w5449_v = ~(v_w5448_v | v_w4769_v);
	assign v_w1093_v = ~(v_w1669_v & v_w1670_v);
	assign v_w3304_v = ~(v_w3126_v & v_w3303_v);
	assign v_w7400_v = ~(v_w1830_v | v_w680_v);
	assign v_w2942_v = ~(v_w2941_v);
	assign v_w3593_v = ~(v_w754_v & v_w2706_v);
	assign v_w72_v = v_s64_v & v_w7107_v;
	assign v_w2591_v = ~(v_w2590_v | v_w617_v);
	assign v_w6668_v = ~(v_w1798_v & v_w1297_v);
	assign v_w3075_v = ~(v_w3072_v | v_w3074_v);
	assign v_w1248_v = ~(v_w8076_v);
	assign v_w6140_v = v_w8062_v ^ v_keyinput_0_v;
	assign v_w6088_v = ~(v_s246_v & v_w889_v);
	assign v_w6635_v = v_w6571_v | v_w1290_v;
	assign v_w6629_v = ~(v_w1188_v | v_w1797_v);
	assign v_w4985_v = ~(v_w4981_v & v_w4984_v);
	assign v_w3504_v = v_w8171_v ^ v_keyinput_75_v;
	assign v_w1928_v = v_s424_v ^ v_w1927_v;
	assign v_w6175_v = v_w6168_v ^ v_w6174_v;
	assign v_w4863_v = ~(v_w555_v & v_w2258_v);
	assign v_w3817_v = ~(v_w2819_v & v_w881_v);
	assign v_w2253_v = ~(v_w2196_v | v_w2191_v);
	assign v_w5787_v = ~(v_s247_v & v_w5786_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s439_v<=0;
	end
	else
	begin
	v_s439_v<=v_w491_v;
	end
	end
	assign v_w223_v = ~(v_w5574_v & v_w5575_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s264_v<=0;
	end
	else
	begin
	v_s264_v<=v_w281_v;
	end
	end
	assign v_w6451_v = ~(v_w6449_v | v_w6450_v);
	assign v_w6064_v = v_w6063_v ^ v_w6033_v;
	assign v_w3969_v = v_w8094_v ^ v_keyinput_22_v;
	assign v_w6617_v = ~(v_w1140_v & v_w1280_v);
	assign v_w1638_v = ~(v_s337_v ^ v_w1154_v);
	assign v_w154_v = v_s145_v & v_w5134_v;
	assign v_w4412_v = ~(v_w1078_v & v_w4411_v);
	assign v_w2978_v = ~(v_s117_v & v_w2355_v);
	assign v_w7154_v = ~(v_w1354_v & v_w7118_v);
	assign v_w55_v = v_s47_v & v_w7107_v;
	assign v_w257_v = ~(v_w7858_v & v_w7859_v);
	assign v_w6193_v = ~(v_w6186_v & v_w6192_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s150_v<=0;
	end
	else
	begin
	v_s150_v<=v_w159_v;
	end
	end
	assign v_w4022_v = ~(v_w4021_v & v_w876_v);
	assign v_w3708_v = ~(v_w3546_v | v_w3707_v);
	assign v_w4132_v = ~(v_w4129_v | v_w4126_v);
	assign v_w7821_v = ~(v_w654_v & v_w7820_v);
	assign v_w7534_v = ~(v_w7265_v & v_w7533_v);
	assign v_w4014_v = ~(v_w3689_v & v_w4010_v);
	assign v_w4159_v = ~(v_w4158_v & v_w690_v);
	assign v_w4151_v = v_s297_v & v_w4054_v;
	assign v_w3113_v = ~(v_w2659_v & v_s387_v);
	assign v_w7414_v = ~(v_w7412_v | v_w7413_v);
	assign v_w3278_v = ~(v_w2541_v ^ v_w2544_v);
	assign v_w6406_v = ~(v_w6399_v | v_w6405_v);
	assign v_w6725_v = ~(v_s412_v & v_w656_v);
	assign v_w3054_v = ~(v_w2358_v & v_s407_v);
	assign v_w5657_v = ~(v_w420_v & v_w3025_v);
	assign v_w5358_v = ~(v_w5126_v & v_w4980_v);
	assign v_w2040_v = ~(v_w2030_v & v_w1100_v);
	assign v_w4569_v = ~(v_w782_v & v_w4568_v);
	assign v_w2283_v = ~(v_s250_v | v_w2268_v);
	assign v_w6010_v = ~(v_w6008_v | v_w6009_v);
	assign v_w1589_v = ~(v_w566_v | v_w578_v);
	assign v_w4774_v = ~(v_w2342_v | v_w4773_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s494_v<=0;
	end
	else
	begin
	v_s494_v<=v_w286_v;
	end
	end
	assign v_w5042_v = ~(v_w5041_v & v_w878_v);
	assign v_w2274_v = ~(v_w926_v & v_w2149_v);
	assign v_w4273_v = ~(v_w4271_v | v_w4272_v);
	assign v_w990_v = ~(v_w2282_v | v_w2283_v);
	assign v_w4200_v = ~(v_s299_v & v_w4169_v);
	assign v_w2751_v = ~(v_s106_v & v_w2355_v);
	assign v_w5862_v = ~(v_w5860_v & v_w5861_v);
	assign v_w5069_v = ~(v_w2391_v | v_w2370_v);
	assign v_w7646_v = ~(v_w657_v | v_w2123_v);
	assign v_w5003_v = ~(v_w5001_v | v_w5002_v);
	assign v_w3333_v = ~(v_w3331_v & v_w3332_v);
	assign v_w1301_v = ~(v_s431_v & v_w562_v);
	assign v_w8132_v = ~(v_w3507_v & v_w4540_v);
	assign v_w2501_v = ~(v_w2416_v | v_w538_v);
	assign v_w7206_v = ~(v_s213_v & v_w7112_v);
	assign v_w1506_v = v_w741_v ^ v_w740_v;
	assign v_w1889_v = ~(v_w1812_v & v_w1888_v);
	assign v_w5409_v = ~(v_w683_v & v_w5408_v);
	assign v_w1486_v = ~(v_w1483_v & v_w1485_v);
	assign v_w543_v = ~(v_w2351_v & v_w991_v);
	assign v_w7281_v = ~(v_w687_v | v_w1362_v);
	assign v_w5461_v = ~(v_w683_v & v_w5460_v);
	assign v_w3596_v = ~(v_w3595_v & v_w873_v);
	assign v_w2412_v = ~(v_w2410_v & v_w2411_v);
	assign v_w8114_v = v_w3518_v | v_w3522_v;
	assign v_w4820_v = ~(v_w2347_v & v_w2766_v);
	assign v_w3983_v = v_w8149_v ^ v_keyinput_59_v;
	assign v_w1209_v = ~(v_w612_v & v_s78_v);
	assign v_w5888_v = ~(v_s321_v & v_w529_v);
	assign v_w6785_v = ~(v_w1075_v | v_w6579_v);
	assign v_w5707_v = ~(v_w2135_v);
	assign v_w4603_v = ~(v_w4601_v & v_w4602_v);
	assign v_w940_v = ~(v_w2697_v | v_w812_v);
	assign v_w7393_v = ~(v_w7391_v | v_w7392_v);
	assign v_w6001_v = ~(v_w5999_v & v_w6000_v);
	assign v_w4300_v = ~(v_w2960_v ^ v_s118_v);
	assign v_w6426_v = ~(v_s160_v & v_w6399_v);
	assign v_w5387_v = ~(v_s351_v & v_w5386_v);
	assign v_w8176_v = v_w5525_v | v_w5526_v;
	assign v_w2609_v = ~(v_w2604_v & v_w2608_v);
	assign v_w1952_v = ~(v_s52_v | v_s51_v);
	assign v_w3082_v = ~(v_w558_v & v_w1124_v);
	assign v_w5349_v = ~(v_w2601_v & v_w2575_v);
	assign v_w8252_v = v_w8251_v ^ v_keyinput_126_v;
	assign v_w5552_v = ~(v_w5550_v & v_w5551_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s349_v<=0;
	end
	else
	begin
	v_s349_v<=v_w385_v;
	end
	end
	assign v_w4976_v = v_w3644_v ^ v_w4541_v;
	assign v_w4630_v = ~(v_w4628_v & v_w4629_v);
	assign v_w6310_v = ~(v_w6018_v | v_w1626_v);
	assign v_w7440_v = ~(v_w680_v | v_w1853_v);
	assign v_w2299_v = ~(v_w2262_v & v_w2298_v);
	assign v_w6536_v = ~(v_w6519_v | v_w6535_v);
	assign v_w7963_v = ~(v_s32_v & v_w2143_v);
	assign v_w255_v = ~(v_w5626_v & v_w5627_v);
	assign v_w1907_v = ~(v_w1807_v | v_w1906_v);
	assign v_w7918_v = ~(v_w527_v & v_w1834_v);
	assign v_w7917_v = ~(v_s87_v & v_w6015_v);
	assign v_w1279_v = ~(v_w874_v & v_s445_v);
	assign v_w1906_v = ~(v_w1904_v & v_w1905_v);
	assign v_w6800_v = v_w656_v & v_s355_v;
	assign v_w2865_v = ~(v_w2862_v & v_w2864_v);
	assign v_w3418_v = ~(v_w3414_v & v_w3417_v);
	assign v_w4298_v = ~(v_w3128_v | v_w4297_v);
	assign v_w7924_v = ~(v_w527_v & v_w944_v);
	assign v_w3623_v = ~(v_w3622_v & v_w2193_v);
	assign v_w1467_v = v_w591_v ^ v_w752_v;
	assign v_w8236_v = v_w8235_v ^ v_keyinput_117_v;
	assign v_w1012_v = ~(v_w564_v & v_s22_v);
	assign v_w2833_v = ~(v_w2819_v);
	assign v_w2706_v = ~(v_w2704_v & v_w2705_v);
	assign v_w6565_v = ~(v_s420_v & v_w666_v);
	assign v_w6349_v = ~(v_w6347_v & v_w6348_v);
	assign v_w5939_v = ~(v_s475_v | v_w461_v);
	assign v_w614_v = ~(v_w612_v | v_w613_v);
	assign v_w7564_v = ~(v_w1548_v | v_w603_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s236_v<=0;
	end
	else
	begin
	v_s236_v<=v_w249_v;
	end
	end
	assign v_w4815_v = ~(v_w4805_v | v_w4528_v);
	assign v_w7417_v = ~(v_w7415_v | v_w7416_v);
	assign v_w5774_v = ~(v_w5772_v & v_w5773_v);
	assign v_w5673_v = ~(v_w4082_v & v_w2671_v);
	assign v_w859_v = ~(v_w1063_v);
	assign v_w5993_v = ~(v_w2091_v ^ v_w2093_v);
	assign v_w3776_v = ~(v_w881_v | v_w1016_v);
	assign v_w957_v = ~(v_w2965_v & v_w2956_v);
	assign v_w7908_v = ~(v_w651_v & v_w7833_v);
	assign v_w8147_v = ~(v_w527_v & v_w1287_v);
	assign v_w646_v = v_w644_v & v_w645_v;
	assign v_w2641_v = ~(v_w2613_v | v_w337_v);
	assign v_w6572_v = ~(v_w1757_v & v_w1140_v);
	assign v_w7019_v = v_w950_v ^ v_w1028_v;
	assign v_w1314_v = ~(v_w1313_v & v_w809_v);
	assign v_w155_v = v_s146_v & v_w5134_v;
	assign v_w2467_v = ~(v_w1131_v | v_w2327_v);
	assign v_w1990_v = v_w680_v | v_w1778_v;
	assign v_w1668_v = ~(v_w1667_v);
	assign v_w677_v = ~(v_s21_v | v_w684_v);
	assign v_w5299_v = ~(v_w2601_v & v_w2417_v);
	assign v_w2480_v = ~(v_w558_v & v_w2399_v);
	assign v_w4984_v = ~(v_w4983_v & v_w866_v);
	assign v_w6826_v = ~(v_w6825_v & v_w1915_v);
	assign v_w6354_v = ~(v_w6322_v | v_w6326_v);
	assign v_w2395_v = ~(v_w2393_v & v_w2394_v);
	assign v_w6437_v = ~(v_w1424_v & v_w6436_v);
	assign v_w1689_v = ~(v_w1417_v | v_w1688_v);
	assign v_w2568_v = v_w2560_v | v_w2565_v;
	assign v_w1982_v = ~(v_w1972_v & v_w1981_v);
	assign v_w3921_v = ~(v_w3919_v & v_w3920_v);
	assign v_w5832_v = ~(v_w5828_v | v_w5831_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s54_v<=0;
	end
	else
	begin
	v_s54_v<=v_w62_v;
	end
	end
	assign v_w5533_v = ~(v_w683_v & v_w5532_v);
	assign v_w4660_v = ~(v_w4512_v ^ v_w3629_v);
	assign v_w7734_v = ~(v_w7732_v & v_w7733_v);
	assign v_w4302_v = ~(v_w4285_v & v_w4288_v);
	assign v_w7213_v = ~(v_w7211_v | v_w7212_v);
	assign v_w2061_v = ~(v_w1418_v & v_w2060_v);
	assign v_w3483_v = ~(v_w3476_v);
	assign v_w2651_v = ~(v_w2650_v | v_w425_v);
	assign v_w1103_v = ~(v_w710_v);
	assign v_w7301_v = v_w7297_v | v_w7300_v;
	assign v_w804_v = ~(v_w806_v | v_w807_v);
	assign v_w3050_v = ~(v_w3048_v | v_w3049_v);
	assign v_w7764_v = ~(v_w7660_v & v_w6829_v);
	assign v_w2744_v = ~(v_w2742_v & v_w2743_v);
	assign v_w6987_v = ~(v_w6982_v | v_w6986_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s191_v<=0;
	end
	else
	begin
	v_s191_v<=v_w204_v;
	end
	end
	assign v_w5152_v = ~(v_w2284_v | v_w1_v);
	assign v_w7854_v = ~(v_s359_v & v_w1993_v);
	assign v_w478_v = ~(v_w4644_v & v_w4654_v);
	assign v_w7530_v = ~(v_w7261_v | v_w7264_v);
	assign v_w2101_v = ~(v_w2099_v & v_w2100_v);
	assign v_w5709_v = ~(v_w892_v & v_w1003_v);
	assign v_w3408_v = ~(v_w3402_v & v_w3407_v);
	assign v_w5611_v = v_w8208_v ^ v_keyinput_100_v;
	assign v_w1699_v = ~(v_w1694_v | v_w1698_v);
	assign v_w3716_v = ~(v_w3690_v & v_w3715_v);
	assign v_w5570_v = ~(v_s221_v & v_w676_v);
	assign v_w2907_v = ~(v_w2361_v | v_w2906_v);
	assign v_w3282_v = ~(v_w3280_v | v_w3281_v);
	assign v_w711_v = v_s310_v | v_s217_v;
	assign v_w5011_v = ~(v_w5006_v | v_w5010_v);
	assign v_w202_v = ~(v_w5524_v & v_w5533_v);
	assign v_w2624_v = ~(v_w2251_v | v_w2599_v);
	assign v_w7031_v = ~(v_w6592_v & v_w831_v);
	assign v_w5519_v = ~(v_w5517_v | v_w5518_v);
	assign v_w1731_v = ~(v_w1728_v & v_w1730_v);
	assign v_w104_v = ~(v_w7157_v & v_w7158_v);
	assign v_w3162_v = ~(v_w3160_v & v_w3161_v);
	assign v_w3289_v = ~(v_s379_v & v_w1_v);
	assign v_w6770_v = ~(v_w6767_v ^ v_w1882_v);
	assign v_w1979_v = ~(v_w1977_v | v_w1978_v);
	assign v_w5773_v = ~(v_w892_v & v_w919_v);
	assign v_w4503_v = ~(v_w4502_v & v_w3633_v);
	assign v_w1405_v = ~(v_w994_v ^ v_w995_v);
	assign v_w3324_v = ~(v_w3322_v & v_w3323_v);
	assign v_w670_v = ~(v_w669_v | v_w667_v);
	assign v_w6953_v = ~(v_w1798_v & v_w1824_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s431_v<=0;
	end
	else
	begin
	v_s431_v<=v_w482_v;
	end
	end
	assign v_w3735_v = ~(v_w3731_v);
	assign v_w7111_v = ~(v_w1144_v & v_w528_v);
	assign v_w5931_v = ~(v_w5929_v & v_w5930_v);
	assign v_w768_v = ~(v_w770_v | v_w771_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s42_v<=0;
	end
	else
	begin
	v_s42_v<=v_w50_v;
	end
	end
	assign v_w2003_v = ~(v_w1363_v | v_w2002_v);
	assign v_w71_v = v_s63_v & v_w7107_v;
	assign v_w5760_v = ~(v_s401_v & v_w529_v);
	assign v_w3038_v = ~(v_w880_v & v_w569_v);
	assign v_w37_v = ~(v_w5608_v & v_w5609_v);
	assign v_w2731_v = ~(v_w699_v & v_s182_v);
	assign v_w2213_v = ~(v_s139_v | v_s138_v);
	assign v_w2975_v = ~(v_w2973_v & v_w2974_v);
	assign v_w3616_v = ~(v_w3484_v | v_w3615_v);
	assign v_w6498_v = ~(v_w6496_v & v_w6497_v);
	assign v_w7210_v = ~(v_s222_v & v_w7113_v);
	assign v_w7628_v = ~(v_w1753_v | v_w7627_v);
	assign v_w3576_v = v_w3573_v | v_w3575_v;
	assign v_w4577_v = ~(v_w3573_v | v_w4576_v);
	assign v_w4722_v = ~(v_w878_v & v_w4569_v);
	assign v_w5738_v = ~(v_s323_v & v_w529_v);
	assign v_w809_v = ~(v_w808_v);
	assign v_w2719_v = ~(v_w2361_v | v_w2718_v);
	assign v_w392_v = ~(v_w6836_v & v_w6850_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s353_v<=0;
	end
	else
	begin
	v_s353_v<=v_w391_v;
	end
	end
	assign v_w2868_v = ~(v_w2355_v & v_s119_v);
	assign v_w4508_v = ~(v_w4450_v & v_w4507_v);
	assign v_w138_v = v_s129_v & v_w5134_v;
	assign v_w2807_v = v_w2806_v ^ v_w553_v;
	assign v_w6810_v = ~(v_w758_v & v_w6804_v);
	assign v_w4054_v = ~(v_w4040_v | v_w885_v);
	assign v_w7707_v = ~(v_w1919_v | v_w7706_v);
	assign v_w7087_v = ~(v_w7083_v | v_w7086_v);
	assign v_w2582_v = ~(v_w2361_v | v_w2581_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s396_v<=0;
	end
	else
	begin
	v_s396_v<=v_w445_v;
	end
	end
	assign v_w2906_v = ~(v_s328_v ^ v_w2643_v);
	assign v_w2128_v = ~(v_w1784_v & v_w2107_v);
	assign v_w2115_v = ~(v_w1783_v & v_w1972_v);
	assign v_w6089_v = ~(v_w657_v & v_s271_v);
	assign v_w2567_v = ~(v_w2547_v & v_w2566_v);
	assign v_w3078_v = ~(v_w558_v & v_w3077_v);
	assign v_w2884_v = ~(v_w2883_v);
	assign v_w7555_v = v_w680_v ^ v_w1378_v;
	assign v_w5147_v = ~(v_w3477_v & v_w5146_v);
	assign v_w2014_v = v_w1026_v & v_w2012_v;
	assign v_w1177_v = ~(v_s85_v | v_s96_v);
	assign v_w2573_v = ~(v_w2570_v | v_w2572_v);
	assign v_w5022_v = ~(v_w5017_v | v_w4589_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s437_v<=0;
	end
	else
	begin
	v_s437_v<=v_w489_v;
	end
	end
	assign v_w225_v = ~(v_w5572_v & v_w5573_v);
	assign v_w1704_v = ~(v_w808_v | v_w1703_v);
	assign v_w5876_v = ~(v_s285_v & v_w528_v);
	assign v_w6823_v = ~(v_w6821_v | v_w6822_v);
	assign v_w8053_v = ~(v_w8007_v | v_w8008_v);
	assign v_w7039_v = ~(v_w1787_v & v_w578_v);
	assign v_w743_v = ~(v_w1102_v & v_w1031_v);
	assign v_w7801_v = ~(v_w6717_v & v_w7800_v);
	assign v_w1769_v = ~(v_w1763_v & v_w1768_v);
	assign v_w3149_v = ~(v_w2860_v ^ v_w2865_v);
	assign v_w3336_v = v_w2497_v ^ v_w2492_v;
	assign v_w644_v = v_w611_v | v_w2028_v;
	assign v_w5919_v = ~(v_w5917_v & v_w5918_v);
	assign v_w4478_v = ~(v_w2910_v | v_w2901_v);
	assign v_w7120_v = v_s20_v & v_w7113_v;
	assign v_w6615_v = ~(v_w6613_v | v_w6614_v);
	assign v_w2323_v = ~(v_w568_v | v_w2322_v);
	assign v_w4982_v = ~(v_w2803_v ^ v_w4400_v);
	assign v_w4402_v = ~(v_w2827_v & v_w4401_v);
	assign v_w1645_v = ~(v_w1374_v | v_w1644_v);
	assign v_w3323_v = ~(v_s313_v & v_w1_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s211_v<=0;
	end
	else
	begin
	v_s211_v<=v_w224_v;
	end
	end
	assign v_w4145_v = ~(v_w2289_v ^ v_s294_v);
	assign v_w4072_v = ~(v_w4070_v & v_w4071_v);
	assign v_w4978_v = ~(v_w2448_v & v_w2585_v);
	assign v_w5343_v = ~(v_w5017_v | v_w5123_v);
	assign v_w8054_v = ~(v_w7981_v | v_w7982_v);
	assign v_w1534_v = ~(v_w1531_v | v_w1533_v);
	assign v_w3586_v = ~(v_w3572_v & v_w3585_v);
	assign v_w7070_v = ~(v_w7069_v & v_w884_v);
	assign v_w5435_v = ~(v_w4776_v);
	assign v_w8199_v = v_w2766_v & v_w697_v;
	assign v_w1340_v = ~(v_w1339_v & v_w809_v);
	assign v_w6286_v = ~(v_w6274_v | v_w6285_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s71_v<=0;
	end
	else
	begin
	v_s71_v<=v_w79_v;
	end
	end
	assign v_w3801_v = ~(v_w3799_v | v_w3800_v);
	assign v_w3540_v = ~(v_w3493_v & v_w3539_v);
	assign v_w7184_v = ~(v_w7117_v | v_w1664_v);
	assign v_w5535_v = ~(v_w5271_v & v_w5037_v);
	assign v_w722_v = ~(v_w786_v | v_w787_v);
	assign v_w4080_v = ~(v_w4078_v & v_w4079_v);
	assign v_w5402_v = ~(v_w683_v & v_w5401_v);
	assign v_w4047_v = ~(v_w4043_v | v_w4046_v);
	assign v_w2292_v = ~(v_w2285_v & v_w2291_v);
	assign v_w3872_v = ~(v_w3870_v | v_w3871_v);
	assign v_w7599_v = ~(v_w1658_v & v_w7598_v);
	assign v_w2311_v = ~(v_w2147_v | v_w531_v);
	assign v_w2919_v = ~(v_w2355_v & v_s352_v);
	assign v_w786_v = ~(v_w1774_v | v_w1995_v);
	assign v_w4967_v = v_w4543_v ^ v_w3645_v;
	assign v_w937_v = ~(v_w3187_v & v_w3188_v);
	assign v_w6510_v = ~(v_w6508_v & v_w6509_v);
	assign v_w1074_v = ~(v_w1705_v & v_w1706_v);
	assign v_w2514_v = ~(v_w2512_v | v_w2513_v);
	assign v_w3794_v = ~(v_w3793_v & v_w2967_v);
	assign v_w3925_v = ~(v_w3798_v | v_w3924_v);
	assign v_w5845_v = ~(v_w5843_v & v_w5844_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s408_v<=0;
	end
	else
	begin
	v_s408_v<=v_w457_v;
	end
	end
	assign v_w6523_v = ~(v_s102_v ^ v_w1700_v);
	assign v_w4004_v = ~(v_w3595_v);
	assign v_w3117_v = ~(v_w699_v & v_s189_v);
	assign v_w1514_v = ~(v_s284_v ^ v_w1513_v);
	assign v_w168_v = ~(v_w7754_v & v_w7755_v);
	assign v_w2238_v = ~(v_s169_v ^ v_w2237_v);
	assign v_w2475_v = v_w2383_v ^ v_w2474_v;
	assign v_w7394_v = v_w7390_v | v_w7393_v;
	assign v_w3146_v = ~(v_w2635_v | v_w3073_v);
	assign v_w7040_v = ~(v_w1798_v & v_w1026_v);
	assign v_w4243_v = ~(v_w4241_v & v_w4242_v);
	assign v_w1002_v = v_w808_v | v_w1288_v;
	assign v_w302_v = ~(v_w7221_v & v_w7222_v);
	assign v_w4137_v = ~(v_w2289_v ^ v_s231_v);
	assign v_w1056_v = ~(v_in11_v ^ v_w1210_v);
	assign v_w1052_v = v_w1051_v;
	assign v_w4060_v = ~(v_w2330_v ^ v_s255_v);
	assign v_w3198_v = ~(v_w3196_v & v_w3197_v);
	assign v_w5468_v = ~(v_w4863_v | v_w4733_v);
	assign v_w7146_v = ~(v_w7118_v & v_w1329_v);
	assign v_w4258_v = ~(v_w3238_v | v_w4257_v);
	assign v_w6038_v = ~(v_w6037_v & v_w6029_v);
	assign v_w5516_v = ~(v_s188_v & v_w5293_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s269_v<=0;
	end
	else
	begin
	v_s269_v<=v_w286_v;
	end
	end
	assign v_w4479_v = ~(v_w4477_v | v_w4478_v);
	assign v_w5155_v = ~(v_w5146_v & v_w1277_v);
	assign v_w3737_v = ~(v_w3734_v | v_w3736_v);
	assign v_w7509_v = ~(v_w679_v & v_w1337_v);
	assign v_w6385_v = ~(v_w6344_v & v_w6343_v);
	assign v_w982_v = ~(v_w1525_v & v_w1526_v);
	assign v_w3934_v = ~(v_w3735_v & v_w3025_v);
	assign v_w6598_v = ~(v_w1751_v & v_w6597_v);
	assign v_w7985_v = ~(v_s469_v | v_s370_v);
	assign v_w927_v = v_s349_v | v_s348_v;
	assign v_w4328_v = ~(v_w3264_v | v_w4327_v);
	assign v_w6238_v = v_s308_v ^ v_w1474_v;
	assign v_w3112_v = ~(v_w3110_v & v_w3111_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s194_v<=0;
	end
	else
	begin
	v_s194_v<=v_w207_v;
	end
	end
	assign v_w4246_v = ~(v_w4245_v & v_w692_v);
	assign v_w1878_v = ~(v_w1876_v & v_w1877_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s275_v<=0;
	end
	else
	begin
	v_s275_v<=v_w293_v;
	end
	end
	assign v_w5000_v = ~(v_w2447_v & v_w2367_v);
	assign v_w1230_v = ~(v_s115_v & v_w1192_v);
	assign v_w2463_v = ~(v_w2461_v | v_w2462_v);
	assign v_w3837_v = ~(v_w2562_v & v_w3732_v);
	assign v_w7946_v = ~(v_w527_v & v_w1435_v);
	assign v_w6690_v = ~(v_w6689_v & v_w655_v);
	assign v_w8117_v = v_w7694_v | v_w7695_v;
	assign v_w7937_v = ~(v_s198_v & v_w2143_v);
	assign v_w4153_v = ~(v_w2554_v);
	assign v_w6022_v = ~(v_s35_v | v_w6021_v);
	assign v_w3134_v = ~(v_w3121_v | v_w1088_v);
	assign v_w2947_v = v_w2940_v | v_w2946_v;
	assign v_w2243_v = ~(v_w2235_v | v_w2242_v);
	assign v_w4009_v = ~(v_w3742_v & v_w4008_v);
	assign v_w3258_v = ~(v_w755_v & v_w2639_v);
	assign v_w5163_v = ~(v_w5146_v & v_w1289_v);
	assign v_w5332_v = ~(v_w2340_v & v_w5037_v);
	assign v_w6961_v = ~(v_w6951_v | v_w6960_v);
	assign v_w3009_v = ~(v_w699_v & v_s180_v);
	assign v_w6869_v = ~(v_w6867_v | v_w6868_v);
	assign v_w3474_v = ~(v_w3472_v & v_w3473_v);
	assign v_w4361_v = ~(v_w4352_v | v_w4360_v);
	assign v_w5265_v = v_s1_v | v_w2332_v;
	assign v_w4783_v = ~(v_w4780_v | v_w4782_v);
	assign v_w4711_v = ~(v_w674_v | v_w4710_v);
	assign v_w7130_v = ~(v_w7128_v | v_w7129_v);
	assign v_w3142_v = ~(v_w3060_v);
	assign v_w4185_v = v_w4181_v ^ v_w4184_v;
	assign v_w4098_v = ~(v_w2312_v & v_w887_v);
	assign v_w4717_v = ~(v_w4715_v & v_w4716_v);
	assign v_w4017_v = ~(v_w4013_v & v_w4016_v);
	assign v_w8187_v = v_w1311_v | v_w6608_v;
	assign v_w6375_v = ~(v_w6374_v & v_w6020_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s182_v<=0;
	end
	else
	begin
	v_s182_v<=v_w195_v;
	end
	end
	assign v_w6894_v = v_w1661_v ^ v_w1659_v;
	assign v_w5757_v = ~(v_w1699_v | v_w5734_v);
	assign v_w3188_v = ~(v_w558_v & v_w3118_v);
	assign v_w5639_v = ~(v_w420_v & v_w2833_v);
	assign v_w4846_v = ~(v_w2369_v & v_w2791_v);
	assign v_w3044_v = ~(v_w3042_v | v_w3043_v);
	assign v_w1631_v = ~(v_s203_v & v_w562_v);
	assign v_w6179_v = ~(v_w664_v & v_s460_v);
	assign v_w2347_v = ~(v_w2261_v);
	assign v_w4590_v = ~(v_w4524_v | v_w4589_v);
	assign v_w1586_v = ~(v_w596_v | v_w602_v);
	assign v_w4108_v = v_s279_v ^ v_w2312_v;
	assign v_w985_v = ~(v_w2021_v | v_w2022_v);
	assign v_w1738_v = ~(v_w1353_v | v_w1737_v);
	assign v_w4683_v = ~(v_w2369_v & v_w2706_v);
	assign v_w1813_v = ~(v_w1373_v);
	assign v_w2909_v = ~(v_w2355_v & v_s200_v);
	assign v_w4385_v = v_w4384_v ^ v_w866_v;
	assign v_w943_v = ~(v_w720_v & v_w942_v);
	assign v_w4234_v = ~(v_w4225_v | v_w4233_v);
	assign v_w4370_v = ~(v_w4367_v & v_w4369_v);
	assign v_w4821_v = ~(v_w4819_v & v_w4820_v);
	assign v_w8213_v = ~(v_w2341_v & v_w673_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s245_v<=0;
	end
	else
	begin
	v_s245_v<=v_w258_v;
	end
	end
	assign v_w1268_v = ~(v_w1266_v & v_w1267_v);
	assign v_w5447_v = ~(v_w5445_v | v_w5446_v);
	assign v_w6219_v = ~(v_s306_v ^ v_w6218_v);
	assign v_o9_v = v_w8168_v ^ v_keyinput_73_v;
	assign v_w3320_v = ~(v_w2619_v | v_w2606_v);
	assign v_w4012_v = ~(v_w4011_v & v_w3689_v);
	assign v_w1895_v = ~(v_w1894_v & v_w1337_v);
	assign v_w5696_v = ~(v_w1496_v | v_w2135_v);
	assign v_w7531_v = ~(v_w7529_v | v_w7530_v);
	assign v_w3274_v = ~(v_w3272_v | v_w3273_v);
	assign v_w5814_v = ~(v_w5812_v & v_w5813_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s499_v<=0;
	end
	else
	begin
	v_s499_v<=v_w336_v;
	end
	end
	assign v_w89_v = ~(v_w7895_v & v_w7896_v);
	assign v_w7551_v = ~(v_w687_v | v_w7239_v);
	assign v_w97_v = ~(v_w7885_v & v_w7886_v);
	assign v_w7500_v = ~(v_w7282_v | v_w7285_v);
	assign v_w4924_v = ~(v_w2369_v & v_w2937_v);
	assign v_w1651_v = ~(v_w1642_v | v_w1650_v);
	assign v_w3915_v = ~(v_w3914_v & v_w957_v);
	assign v_w7252_v = ~(v_w7250_v | v_w7251_v);
	assign v_w5180_v = ~(v_w693_v | v_w2238_v);
	assign v_w6079_v = ~(v_s359_v & v_w6050_v);
	assign v_w4541_v = ~(v_w8133_v);
	assign v_o21_v = ~(v_s219_v ^ v_s2_v);
	assign v_w4411_v = ~(v_w1079_v | v_w4410_v);
	assign v_w1520_v = ~(v_w1518_v & v_w1519_v);
	assign v_w7277_v = ~(v_w680_v & v_w1066_v);
	assign v_w2005_v = ~(v_w2004_v | v_w1725_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s365_v<=0;
	end
	else
	begin
	v_s365_v<=v_w408_v;
	end
	end
	assign v_w3091_v = ~(v_w3089_v & v_w3090_v);
	assign v_w7399_v = ~(v_w687_v | v_w566_v);
	assign v_w7312_v = ~(v_w679_v | v_w895_v);
	assign v_w3813_v = ~(v_w2856_v | v_w881_v);
	assign v_w6100_v = ~(v_w6099_v ^ v_s273_v);
	assign v_w301_v = ~(v_w5628_v & v_w5629_v);
	assign v_w7887_v = ~(v_s109_v & v_w7876_v);
	assign v_w3547_v = ~(v_w3546_v);
	assign v_w7323_v = ~(v_w679_v | v_w1401_v);
	assign v_w4983_v = ~(v_w4863_v | v_w4982_v);
	assign v_w6030_v = ~(v_w657_v | v_w396_v);
	assign v_w7916_v = ~(v_w527_v & v_w607_v);
	assign v_w6724_v = ~(v_w6722_v | v_w6723_v);
	assign v_w1815_v = ~(v_w1699_v & v_w1075_v);
	assign v_w198_v = ~(v_w5480_v & v_w5487_v);
	assign v_w514_v = ~(v_w6222_v & v_w6232_v);
	assign v_w3758_v = v_w2706_v | v_w3735_v;
	assign v_w2205_v = ~(v_s149_v | v_s148_v);
	assign v_w5363_v = ~(v_w4965_v & v_w5126_v);
	assign v_w7413_v = ~(v_w575_v | v_w680_v);
	assign v_w5950_v = ~(v_w5707_v & v_w1638_v);
	assign v_w1360_v = ~(v_w1356_v | v_w1359_v);
	assign v_w5836_v = ~(v_w2117_v & v_w1021_v);
	assign v_w7375_v = ~(v_w7373_v | v_w7374_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s489_v<=0;
	end
	else
	begin
	v_s489_v<=v_w184_v;
	end
	end
	assign v_w129_v = ~(v_w5646_v & v_w5647_v);
	assign v_w6969_v = v_w1598_v ^ v_w6962_v;
	assign v_w6144_v = ~(v_w6142_v & v_w6143_v);
	assign v_w406_v = ~(v_w4284_v & v_w4290_v);
	assign v_w6133_v = ~(v_s244_v & v_w6105_v);
	assign v_w659_v = ~(v_w657_v | v_w658_v);
	assign v_w267_v = ~(v_w5305_v & v_w5313_v);
	assign v_w515_v = ~(v_w6248_v & v_w6259_v);
	assign v_w7090_v = ~(v_w7087_v & v_w7089_v);
	assign v_w5525_v = ~(v_w3199_v | v_w2370_v);
	assign v_w2619_v = ~(v_w2618_v);
	assign v_w6228_v = ~(v_w6198_v | v_w6227_v);
	assign v_w5812_v = ~(v_w5811_v & v_w2113_v);
	assign v_w7102_v = ~(v_w5906_v | v_w7101_v);
	assign v_w6798_v = ~(v_w6797_v & v_w655_v);
	assign v_w577_v = ~(v_w665_v & v_s243_v);
	assign v_w825_v = ~(v_w823_v | v_w824_v);
	assign v_w4142_v = ~(v_w887_v & v_w2290_v);
	assign v_w6149_v = ~(v_w6147_v | v_w6148_v);
	assign v_w5177_v = v_w5141_v & v_s76_v;
	assign v_w6265_v = ~(v_w6264_v & v_w6020_v);
	assign v_w116_v = ~(v_w7772_v & v_w7773_v);
	assign v_w3065_v = ~(v_w2484_v & v_w3060_v);
	assign v_w3835_v = ~(v_w3833_v & v_w3834_v);
	assign v_w2870_v = v_s360_v ^ v_w2645_v;
	assign v_w5669_v = ~(v_w420_v & v_w2706_v);
	assign v_w6087_v = ~(v_w6085_v | v_w6086_v);
	assign v_w3087_v = ~(v_w3085_v | v_w3086_v);
	assign v_w3954_v = ~(v_w3952_v | v_w3953_v);
	assign v_w6951_v = ~(v_w6949_v & v_w6950_v);
	assign v_w6008_v = ~(v_w6006_v & v_w6007_v);
	assign v_w6648_v = ~(v_w6647_v & v_w6626_v);
	assign v_w1910_v = ~(v_w1187_v | v_w893_v);
	assign v_w5550_v = ~(v_w4431_v | v_w5549_v);
	assign v_w5161_v = v_w5141_v & v_s22_v;
	assign v_w1352_v = ~(v_w1342_v & v_w1351_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s280_v<=0;
	end
	else
	begin
	v_s280_v<=v_w299_v;
	end
	end
	assign v_w1551_v = ~(v_w1549_v & v_w1550_v);
	assign v_w1240_v = ~(v_s346_v & v_w1103_v);
	assign v_w4359_v = ~(v_w690_v & v_w4358_v);
	assign v_w6449_v = ~(v_w5999_v & v_w6448_v);
	assign v_w4441_v = ~(v_w4439_v & v_w4440_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s256_v<=0;
	end
	else
	begin
	v_s256_v<=v_w271_v;
	end
	end
	assign v_w7445_v = ~(v_w7443_v | v_w7444_v);
	assign v_w1880_v = ~(v_w1878_v & v_w1879_v);
	assign v_w5703_v = v_w2113_v;
	assign v_w5379_v = ~(v_w4863_v | v_w4933_v);
	assign v_w5668_v = ~(v_s423_v & v_w695_v);
	assign v_w5972_v = ~(v_w892_v & v_w1074_v);
	assign v_w3555_v = ~(v_w3551_v & v_w3554_v);
	assign v_w5414_v = ~(v_w4848_v | v_w5123_v);
	assign v_w8188_v = v_w758_v ^ v_keyinput_88_v;
	assign v_w791_v = ~(v_w2167_v & v_w2173_v);
	assign v_w3356_v = ~(v_w3354_v | v_w3355_v);
	assign v_w871_v = ~(v_w1012_v & v_w1013_v);
	assign v_w2657_v = ~(v_w2656_v | v_w432_v);
	assign v_w965_v = ~(v_w3189_v & v_w3190_v);
	assign v_w2235_v = ~(v_w2234_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s447_v<=0;
	end
	else
	begin
	v_s447_v<=v_w500_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s261_v<=0;
	end
	else
	begin
	v_s261_v<=v_w277_v;
	end
	end
	assign v_w5025_v = ~(v_w5023_v & v_w5024_v);
	assign v_w2455_v = ~(v_w2242_v | v_w2234_v);
	assign v_w2096_v = ~(v_w2094_v | v_w2095_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s127_v<=0;
	end
	else
	begin
	v_s127_v<=v_w136_v;
	end
	end
	assign v_w1319_v = ~(v_w875_v & v_s437_v);
	assign v_w528_v = ~(v_s475_v);
	assign v_w2006_v = v_w1725_v & v_w2004_v;
	assign v_w5587_v = ~(v_w675_v & v_w5416_v);
	assign v_w1614_v = ~(v_w953_v & v_w1613_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s2_v<=0;
	end
	else
	begin
	v_s2_v<=v_w2_v;
	end
	end
	assign v_w7297_v = ~(v_w7295_v | v_w7296_v);
	assign v_w7855_v = ~(v_w651_v & v_w7672_v);
	assign v_w8012_v = ~(v_w8010_v & v_w8011_v);
	assign v_w5544_v = ~(v_w4431_v | v_w5543_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s27_v<=0;
	end
	else
	begin
	v_s27_v<=v_w30_v;
	end
	end
	assign v_w380_v = ~(v_w6887_v & v_w6888_v);
	assign v_w855_v = ~(v_w853_v | v_w854_v);
	assign v_w617_v = ~(v_w605_v & v_w556_v);
	assign v_w7038_v = ~(v_w6602_v | v_w7037_v);
	assign v_w3641_v = ~(v_w3491_v | v_w3537_v);
	assign v_w3181_v = ~(v_w3176_v | v_w3180_v);
	assign v_w345_v = ~(v_s500_v);
	assign v_w6261_v = ~(v_w6238_v & v_w6237_v);
	assign v_w6431_v = ~(v_w6430_v & v_w659_v);
	assign v_w1548_v = v_w567_v ^ v_w578_v;
	assign v_w621_v = ~(v_w2725_v | v_w2728_v);
	assign v_w3792_v = ~(v_w3787_v & v_w3790_v);
	assign v_w3256_v = ~(v_w2635_v | v_w2686_v);
	assign v_w7319_v = ~(v_w679_v | v_w847_v);
	assign v_w7283_v = ~(v_w687_v | v_w1729_v);
	assign v_w2180_v = ~(v_w2165_v | v_w2179_v);
	assign v_w6441_v = ~(v_w6029_v | v_w6440_v);
	assign v_w5151_v = ~(v_w8101_v);
	assign v_w6138_v = ~(v_w6124_v | v_w6137_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s11_v<=0;
	end
	else
	begin
	v_s11_v<=v_w12_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s147_v<=0;
	end
	else
	begin
	v_s147_v<=v_w156_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s281_v<=0;
	end
	else
	begin
	v_s281_v<=v_w300_v;
	end
	end
	assign v_w6212_v = v_w1490_v ^ v_w6211_v;
	assign v_w6984_v = ~(v_w6983_v & v_w1915_v);
	assign v_w5061_v = ~(v_w5059_v | v_w5060_v);
	assign v_w8116_v = v_w8115_v ^ v_keyinput_38_v;
	assign v_w2989_v = v_w552_v ^ v_w2988_v;
	assign v_w974_v = ~(v_w1024_v | v_w978_v);
	assign v_w599_v = ~(v_w597_v | v_w598_v);
	assign v_w237_v = ~(v_w7866_v & v_w7867_v);
	assign v_w7411_v = ~(v_w7406_v & v_w7409_v);
	assign v_w7215_v = ~(v_w1514_v | v_w528_v);
	assign v_w5254_v = ~(v_w8116_v);
	assign v_w7117_v = ~(v_w528_v & v_w612_v);
	assign v_w516_v = ~(v_w6265_v & v_w6286_v);
	assign v_w4850_v = ~(v_w4847_v | v_w4849_v);
	assign v_w6207_v = ~(v_w664_v & v_s461_v);
	assign v_w340_v = ~(v_w4198_v & v_w4204_v);
	assign v_w636_v = v_w639_v & v_w640_v;
	assign v_w3686_v = ~(v_w3451_v & v_w3483_v);
	assign v_w416_v = ~(v_w4328_v & v_w4345_v);
	assign v_w2715_v = ~(v_w699_v & v_s183_v);
	assign v_w3671_v = ~(v_w3632_v & v_w3670_v);
	assign v_w2411_v = ~(v_w698_v & v_s254_v);
	assign v_w2281_v = ~(v_w2279_v | v_w2280_v);
	assign v_w744_v = v_in31_v ^ v_w777_v;
	assign v_w3445_v = ~(v_w3443_v & v_w3444_v);
	assign v_w2603_v = ~(v_w2596_v & v_w1139_v);
	assign v_w4464_v = ~(v_w2558_v | v_w2367_v);
	assign v_w5218_v = ~(v_w5216_v | v_w5217_v);
	assign v_w6971_v = ~(v_w6968_v | v_w6970_v);
	assign v_w1088_v = ~(v_w1086_v | v_w1087_v);
	assign v_w3036_v = ~(v_w3035_v | v_w557_v);
	assign v_w3024_v = ~(v_w558_v & v_w1079_v);
	assign v_w2371_v = ~(v_w2368_v | v_w2370_v);
	assign v_w3165_v = ~(v_w3163_v & v_w3164_v);
	assign v_w6408_v = ~(v_w6406_v | v_w6407_v);
	assign v_w4684_v = ~(v_w4682_v & v_w4683_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s93_v<=0;
	end
	else
	begin
	v_s93_v<=v_w101_v;
	end
	end
	assign v_w5716_v = ~(v_w5712_v | v_w5715_v);
	assign v_w1031_v = ~(v_w1029_v & v_w1030_v);
	assign v_w5489_v = ~(v_w4655_v);
	assign v_w5127_v = ~(v_w878_v | v_w5126_v);
	assign v_w2985_v = ~(v_w2984_v);
	assign v_w280_v = ~(v_s493_v);
	assign v_w2322_v = ~(v_w2321_v);
	assign v_w3290_v = ~(v_w3288_v & v_w3289_v);
	assign v_w6925_v = ~(v_w6923_v | v_w6924_v);
	assign v_w1123_v = ~(v_w2300_v & v_w1329_v);
	assign v_w3700_v = ~(v_w3694_v | v_w3699_v);
	assign v_w479_v = ~(v_w4598_v & v_w4615_v);
	assign v_w2778_v = ~(v_w2148_v & v_w2777_v);
	assign v_w1329_v = ~(v_w770_v ^ v_w771_v);
	assign v_o10_v = v_w8033_v ^ v_w8061_v;
	assign v_w7999_v = ~(v_s461_v | v_s311_v);
	assign v_w7780_v = ~(v_w6768_v | v_w1919_v);
	assign v_w1781_v = ~(v_w685_v);
	assign v_w2380_v = ~(v_w2379_v | v_w2296_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s383_v<=0;
	end
	else
	begin
	v_s383_v<=v_w429_v;
	end
	end
	assign v_w3157_v = ~(v_w3121_v | v_w2856_v);
	assign v_w669_v = ~(v_w730_v);
	assign v_w1119_v = ~(v_w1117_v & v_w1118_v);
	assign v_w6799_v = ~(v_w1397_v | v_w6571_v);
	assign v_w3846_v = ~(v_w2308_v & v_w3732_v);
	assign v_w1840_v = ~(v_w1833_v | v_w1839_v);
	assign v_w3610_v = ~(v_w3199_v | v_w1068_v);
	assign v_w6673_v = ~(v_w656_v & v_s437_v);
	assign v_w6448_v = ~(v_w664_v & v_s469_v);
	assign v_w234_v = ~(v_w5570_v & v_w5571_v);
	assign v_w676_v = ~(v_w675_v);
	assign v_w233_v = ~(v_w5347_v & v_w5353_v);
	assign v_w4146_v = ~(v_s281_v & v_w4116_v);
	assign v_w799_v = v_w797_v | v_w798_v;
	assign v_w633_v = v_w1126_v & v_w2054_v;
	assign v_w2633_v = ~(v_w2629_v & v_w2632_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s126_v<=0;
	end
	else
	begin
	v_s126_v<=v_w135_v;
	end
	end
	assign v_w4888_v = v_w3643_v ^ v_w4482_v;
	assign v_w5370_v = ~(v_s201_v & v_w5293_v);
	assign v_w7795_v = ~(v_w7793_v & v_w7794_v);
	assign v_w1451_v = ~(v_w1447_v | v_w1450_v);
	assign v_w4870_v = ~(v_w4869_v & v_w878_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s153_v<=0;
	end
	else
	begin
	v_s153_v<=v_w162_v;
	end
	end
	assign v_w7163_v = ~(v_w1701_v | v_w529_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s128_v<=0;
	end
	else
	begin
	v_s128_v<=v_w137_v;
	end
	end
	assign v_w158_v = v_s149_v & v_w5134_v;
	assign v_w197_v = ~(v_w5472_v & v_w5479_v);
	assign v_w5539_v = ~(v_w5537_v | v_w5538_v);
	assign v_w5159_v = ~(v_w1136_v & v_s1_v);
	assign v_w6793_v = ~(v_w1816_v | v_w6608_v);
	assign v_w6923_v = ~(v_w6602_v | v_w6922_v);
	assign v_w7641_v = v_w7640_v ^ v_w1378_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s330_v<=0;
	end
	else
	begin
	v_s330_v<=v_w358_v;
	end
	end
	assign v_w8189_v = ~(v_w596_v | v_w1782_v);
	assign v_w5851_v = ~(v_w5849_v | v_w5850_v);
	assign v_w2734_v = ~(v_s381_v ^ v_w2652_v);
	assign v_w1269_v = ~(v_s274_v & v_w1192_v);
	assign v_w951_v = ~(v_w1487_v & v_w1598_v);
	assign v_w3424_v = ~(v_w2607_v & v_w2690_v);
	assign v_w6416_v = ~(v_w6414_v & v_w6415_v);
	assign v_w1916_v = ~(v_w1912_v & v_w1915_v);
	assign v_w7129_v = ~(v_w528_v | v_w888_v);
	assign v_w6121_v = ~(v_w5746_v & v_w6120_v);
	assign v_w6571_v = ~(v_w1972_v & v_w1986_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s293_v<=0;
	end
	else
	begin
	v_s293_v<=v_w315_v;
	end
	end
	assign v_w3663_v = ~(v_w3641_v & v_w3662_v);
	assign v_w7781_v = ~(v_w1883_v | v_w1782_v);
	assign v_w4805_v = v_w4534_v ^ v_w4494_v;
	assign v_w6541_v = ~(v_w6539_v & v_w6540_v);
	assign v_w6102_v = ~(v_s246_v & v_w1557_v);
	assign v_w5144_v = ~(v_w5142_v | v_w5143_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s108_v<=0;
	end
	else
	begin
	v_s108_v<=v_w116_v;
	end
	end
	assign v_w6880_v = ~(v_w6876_v | v_w6879_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s177_v<=0;
	end
	else
	begin
	v_s177_v<=v_w190_v;
	end
	end
	assign v_w3747_v = ~(v_w964_v | v_w3735_v);
	assign v_w3041_v = v_w3040_v ^ v_w553_v;
	assign v_w5662_v = ~(v_s84_v & v_w695_v);
	assign v_w4900_v = ~(v_w4898_v | v_w4899_v);
	assign v_w1644_v = ~(v_s334_v ^ v_w1643_v);
	assign v_w7617_v = ~(v_w7615_v | v_w7616_v);
	assign v_w2891_v = ~(v_w2484_v & v_w2890_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s277_v<=0;
	end
	else
	begin
	v_s277_v<=v_w296_v;
	end
	end
	assign v_w3675_v = ~(v_w1008_v & v_w3674_v);
	assign v_w7835_v = ~(v_s446_v & v_w7742_v);
	assign v_w4495_v = ~(v_w4455_v & v_w4494_v);
	assign v_w1927_v = ~(v_w780_v & v_s7_v);
	assign v_w7360_v = ~(v_w7358_v | v_w7359_v);
	assign v_w2389_v = ~(v_w699_v & v_s238_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s289_v<=0;
	end
	else
	begin
	v_s289_v<=v_w309_v;
	end
	end
	assign v_w4197_v = ~(v_w2799_v | v_w4041_v);
	assign v_w7140_v = ~(v_w528_v | v_w1928_v);
	assign v_w998_v = ~(v_w997_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s415_v<=0;
	end
	else
	begin
	v_s415_v<=v_w466_v;
	end
	end
	assign v_w2179_v = ~(v_s170_v | v_w2178_v);
	assign v_w1684_v = ~(v_w1094_v | v_w1678_v);
	assign v_w3806_v = ~(v_w572_v | v_w3735_v);
	assign v_w2635_v = ~(v_w2634_v);
	assign v_w5153_v = v_w5140_v & v_s14_v;
	assign v_w7173_v = ~(v_w7171_v | v_w7172_v);
	assign v_w1135_v = ~(v_w1134_v);
	assign v_w7024_v = ~(v_w7020_v | v_w7023_v);
	assign v_w3654_v = ~(v_w3651_v | v_w3653_v);
	assign v_w4109_v = ~(v_w2321_v & v_s266_v);
	assign v_w7698_v = ~(v_w654_v & v_w7697_v);
	assign v_w4554_v = ~(v_w958_v & v_w4553_v);
	assign v_w4371_v = ~(v_w3017_v ^ v_s391_v);
	assign v_w6905_v = ~(v_w6895_v | v_w6904_v);
	assign v_w3440_v = ~(v_w3438_v | v_w3439_v);
	assign v_w5269_v = ~(v_w1069_v | v_w2264_v);
	assign v_w67_v = v_s59_v & v_w7107_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s515_v<=0;
	end
	else
	begin
	v_s515_v<=v_w436_v;
	end
	end
	assign v_w4039_v = v_w1_v & v_s156_v;
	assign v_w2569_v = ~(v_w2567_v & v_w2568_v);
	assign v_w6753_v = ~(v_w6751_v & v_w6752_v);
	assign v_w6582_v = ~(v_w656_v & v_s451_v);
	assign v_w2840_v = v_w355_v ^ v_w2642_v;
	assign v_w4333_v = ~(v_w4331_v & v_w4332_v);
	assign v_w3436_v = ~(v_w2995_v ^ v_w2996_v);
	assign v_w7819_v = ~(v_w7817_v | v_w7818_v);
	assign v_w5002_v = ~(v_w2619_v | v_w2370_v);
	assign v_w6214_v = ~(v_w6213_v & v_w659_v);
	assign v_w7982_v = v_s471_v & v_s390_v;
	assign v_w2451_v = ~(v_w2371_v | v_w2450_v);
	assign v_w3125_v = ~(v_w1139_v);
	assign v_w2133_v = ~(v_w2132_v | v_w2121_v);
	assign v_w1696_v = ~(v_s399_v ^ v_w1161_v);
	assign v_w8154_v = v_w5279_v | v_w5285_v;
	assign v_w6780_v = ~(v_w6778_v | v_w6779_v);
	assign v_w5028_v = ~(v_w5027_v & v_w673_v);
	assign v_w2674_v = ~(v_w2484_v & v_w2671_v);
	assign v_w4745_v = ~(v_w4744_v & v_w878_v);
	assign v_w4946_v = ~(v_w878_v & v_w4546_v);
	assign v_w5769_v = ~(v_w1101_v | v_w5734_v);
	assign v_w6152_v = ~(v_s286_v & v_w1528_v);
	assign v_w1951_v = ~(v_s54_v | v_s53_v);
	assign v_w2553_v = v_w531_v & v_s291_v;
	assign v_w3106_v = ~(v_w3104_v & v_w3105_v);
	assign v_w4100_v = ~(v_s280_v & v_w4056_v);
	assign v_w4038_v = ~(v_s1_v | v_s40_v);
	assign v_w3975_v = ~(v_w3732_v & v_w3077_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s509_v<=0;
	end
	else
	begin
	v_s509_v<=v_w395_v;
	end
	end
	assign v_w6409_v = ~(v_w1667_v & v_w6378_v);
	assign v_w7836_v = ~(v_w6599_v | v_w1919_v);
	assign v_w5086_v = v_w5085_v & v_w4588_v;
	assign v_w6945_v = v_w656_v & v_s322_v;
	assign v_w2161_v = v_w531_v | v_w2160_v;
	assign v_w5712_v = ~(v_s475_v | v_w373_v);
	assign v_w446_v = ~(v_w4740_v & v_w4755_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s22_v<=0;
	end
	else
	begin
	v_s22_v<=v_w24_v;
	end
	end
	assign v_w1345_v = ~(v_w874_v & v_s412_v);
	assign v_w5820_v = ~(v_w1902_v | v_w2138_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s514_v<=0;
	end
	else
	begin
	v_s514_v<=v_w431_v;
	end
	end
	assign v_o11_v = ~(v_w8030_v ^ v_w8031_v);
	assign v_w7107_v = ~(v_w1972_v & v_w1933_v);
	assign v_w6289_v = ~(v_w6287_v & v_w6288_v);
	assign v_w7723_v = ~(v_w654_v & v_w7722_v);
	assign v_w4097_v = ~(v_w4088_v | v_w4096_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s462_v<=0;
	end
	else
	begin
	v_s462_v<=v_w515_v;
	end
	end
	assign v_w3167_v = v_w2522_v ^ v_w2523_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s250_v<=0;
	end
	else
	begin
	v_s250_v<=v_w264_v;
	end
	end
	assign v_w4928_v = ~(v_w4925_v | v_w4927_v);
	assign v_w2147_v = v_w263_v & v_w946_v;
	assign v_w6353_v = ~(v_w1644_v | v_w6325_v);
	assign v_w2991_v = ~(v_w1083_v);
	assign v_w384_v = ~(v_s507_v);
	assign v_w4963_v = ~(v_w2342_v | v_w4962_v);
	assign v_w1822_v = ~(v_w1095_v & v_w1126_v);
	assign v_w4248_v = ~(v_w3379_v & v_w4247_v);
	assign v_w6603_v = ~(v_w2102_v ^ v_w1908_v);
	assign v_w1305_v = ~(v_w1052_v & v_s26_v);
	assign v_w2009_v = ~(v_w2008_v | v_w1678_v);
	assign v_w4051_v = ~(v_w4050_v | v_s172_v);
	assign v_w3475_v = v_w2358_v & v_s426_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s343_v<=0;
	end
	else
	begin
	v_s343_v<=v_w378_v;
	end
	end
	assign v_w7650_v = ~(v_w7648_v | v_w7649_v);
	assign v_w7524_v = ~(v_w7522_v | v_w7523_v);
	assign v_w8149_v = ~(v_w3981_v & v_w3982_v);
	assign v_w6258_v = ~(v_w6018_v | v_w1474_v);
	assign v_w5327_v = ~(v_w5046_v & v_w5326_v);
	assign v_w6057_v = ~(v_w6056_v & v_w6020_v);
	assign v_w1118_v = ~(v_w562_v & v_s84_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s10_v<=0;
	end
	else
	begin
	v_s10_v<=v_w11_v;
	end
	end
	assign v_w31_v = ~(v_w5610_v & v_w5611_v);
	assign v_w8088_v = v_w3128_v | v_w3131_v;
	assign v_w61_v = v_s53_v & v_w7107_v;
	assign v_w6339_v = ~(v_w6334_v & v_w6338_v);
	assign v_w2442_v = ~(v_w2441_v);
	assign v_w5786_v = ~(v_s475_v & v_w2135_v);
	assign v_w6410_v = ~(v_w6381_v & v_w6379_v);
	assign v_w2124_v = ~(v_w2105_v | v_w2123_v);
	assign v_w1399_v = ~(v_w1396_v | v_w1398_v);
	assign v_w7320_v = ~(v_w1816_v | v_w680_v);
	assign v_w6694_v = v_w1742_v ^ v_w1891_v;
	assign v_w6535_v = ~(v_w6525_v & v_w6534_v);
	assign v_w2472_v = ~(v_w2441_v | v_w2471_v);
	assign v_w4618_v = ~(v_w2667_v | v_w2261_v);
	assign v_w5366_v = ~(v_w4863_v | v_w4962_v);
	assign v_w3302_v = ~(v_w2713_v | v_w762_v);
	assign v_w5685_v = ~(v_w5684_v & v_w2120_v);
	assign v_w4700_v = v_w3631_v ^ v_w4570_v;
	assign v_w3285_v = ~(v_w2346_v & v_w2634_v);
	assign v_w4641_v = ~(v_w4639_v & v_w4640_v);
	assign v_w5223_v = ~(v_s198_v & v_w5140_v);
	assign v_w6661_v = ~(v_w8201_v);
	assign v_w418_v = ~(v_w7173_v & v_w7174_v);
	assign v_w7496_v = ~(v_w7310_v & v_w7495_v);
	assign v_w1158_v = ~(v_w1157_v & v_w373_v);
	assign v_w1789_v = ~(v_w1788_v & v_w1187_v);
	assign v_w5107_v = ~(v_w4588_v & v_w5106_v);
	assign v_w200_v = ~(v_w5508_v & v_w5515_v);
	assign v_w2002_v = ~(v_w1119_v ^ v_w1999_v);
	assign v_w5179_v = ~(v_w5146_v & v_w1339_v);
	assign v_w7651_v = ~(v_w7645_v | v_w7650_v);
	assign v_w313_v = ~(v_w3420_v & v_w3423_v);
	assign v_w6729_v = ~(v_w1886_v ^ v_w1887_v);
	assign v_w6389_v = v_w8162_v ^ v_keyinput_68_v;
	assign v_w244_v = ~(v_w5566_v & v_w5567_v);
	assign v_w2710_v = ~(v_w558_v & v_w753_v);
	assign v_w2928_v = ~(v_s346_v & v_w565_v);
	assign v_w2341_v = ~(v_w2234_v | v_w2257_v);
	assign v_w6056_v = ~(v_s86_v ^ v_w6055_v);
	assign v_w2626_v = ~(v_w2243_v | v_w2625_v);
	assign v_w5695_v = ~(v_w5693_v | v_w5694_v);
	assign v_w896_v = v_w894_v | v_w895_v;
	assign v_w1083_v = ~(v_w1081_v | v_w1082_v);
	assign v_w51_v = ~(v_w5666_v & v_w5667_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s352_v<=0;
	end
	else
	begin
	v_s352_v<=v_w390_v;
	end
	end
	assign v_w7002_v = ~(v_w1788_v & v_w1026_v);
	assign v_w7282_v = ~(v_w8211_v);
	assign v_w7625_v = ~(v_w7624_v & v_w1298_v);
	assign v_w1475_v = ~(v_w1374_v | v_w1474_v);
	assign v_w2008_v = ~(v_w723_v ^ v_w1094_v);
	assign v_w6046_v = ~(v_w6044_v & v_w6045_v);
	assign v_w3692_v = ~(v_w3538_v);
	assign v_w3_v = ~(v_w7913_v & v_w7914_v);
	assign v_w3236_v = ~(v_w2635_v | v_w2718_v);
	assign v_w6778_v = ~(v_w656_v | v_w6777_v);
	assign v_w2498_v = ~(v_w2492_v & v_w2497_v);
	assign v_w5247_v = ~(v_s289_v & v_w5141_v);
	assign v_w485_v = ~(v_w7653_v & v_w7654_v);
	assign v_w4565_v = ~(v_w4563_v | v_w4564_v);
	assign v_w6718_v = ~(v_w884_v & v_w6714_v);
	assign v_w2273_v = ~(v_w2145_v & v_w2152_v);
	assign v_w1477_v = ~(v_w1476_v | v_w808_v);
	assign v_w7833_v = ~(v_w7831_v & v_w7832_v);
	assign v_w102_v = ~(v_w5596_v & v_w5597_v);
	assign v_w4894_v = ~(v_w2956_v | v_w2370_v);
	assign v_w303_v = ~(v_w7217_v & v_w7218_v);
	assign v_w7480_v = ~(v_w7332_v & v_w7329_v);
	assign v_w6118_v = v_w6113_v ^ v_w6117_v;
	assign v_w7219_v = ~(v_w1528_v | v_w528_v);
	assign v_w3015_v = ~(v_s111_v | v_w844_v);
	assign v_w3141_v = ~(v_w3139_v & v_w3140_v);
	assign v_w911_v = ~(v_w2139_v | v_w2142_v);
	assign v_w1449_v = ~(v_w666_v & v_s159_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s123_v<=0;
	end
	else
	begin
	v_s123_v<=v_w132_v;
	end
	end
	assign v_w5008_v = ~(v_w2458_v & v_w5007_v);
	assign v_w8221_v = v_w6864_v | v_w6865_v;
	assign v_w7110_v = ~(v_s7_v & v_w7109_v);
	assign v_w5122_v = ~(v_w5119_v | v_w5121_v);
	assign v_w4838_v = ~(v_w674_v & v_s369_v);
	assign v_w1522_v = ~(v_w1521_v | v_w1180_v);
	assign v_w7922_v = ~(v_w527_v & v_w578_v);
	assign v_w389_v = ~(v_w5387_v & v_w5394_v);
	assign v_w4980_v = ~(v_w3644_v ^ v_w4468_v);
	assign v_w246_v = ~(v_w7698_v & v_w7699_v);
	assign v_w807_v = ~(v_in7_v ^ v_w1198_v);
	assign v_w8228_v = ~(v_w662_v & v_w1337_v);
	assign v_w2803_v = ~(v_w2801_v & v_w2802_v);
	assign v_w6364_v = ~(v_w664_v & v_s466_v);
	assign v_w6312_v = ~(v_w6307_v & v_w6311_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s443_v<=0;
	end
	else
	begin
	v_s443_v<=v_w495_v;
	end
	end
	assign v_w4260_v = ~(v_w2896_v | v_s331_v);
	assign v_w3935_v = ~(v_w3933_v & v_w3934_v);
	assign v_w427_v = ~(v_w3344_v & v_w3351_v);
	assign v_w4392_v = ~(v_w8064_v);
	assign v_w6048_v = ~(v_w396_v | v_s477_v);
	assign v_w6671_v = ~(v_w6662_v & v_w6670_v);
	assign v_w5675_v = ~(v_w4082_v & v_w3100_v);
	assign v_w6732_v = ~(v_w1798_v & v_w1350_v);
	assign v_w1495_v = ~(v_w1493_v & v_w1494_v);
	assign v_w6787_v = ~(v_w1691_v ^ v_w1709_v);
	assign v_w862_v = ~(v_w3014_v & v_w3019_v);
	assign v_w981_v = v_w2027_v & v_w945_v;
	assign v_w6279_v = ~(v_s207_v ^ v_w6278_v);
	assign v_w2210_v = v_w2208_v & v_w2209_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s344_v<=0;
	end
	else
	begin
	v_s344_v<=v_w379_v;
	end
	end
	assign v_w3032_v = ~(v_w3031_v & v_w697_v);
	assign v_w6839_v = ~(v_w1787_v & v_w1453_v);
	assign v_w7454_v = ~(v_w7446_v | v_w7453_v);
	assign v_w5255_v = ~(v_s274_v & v_w5140_v);
	assign v_w2386_v = ~(v_s239_v & v_w2355_v);
	assign v_w7499_v = ~(v_w7301_v & v_w7498_v);
	assign v_w2388_v = ~(v_w2358_v & v_s281_v);
	assign v_w7479_v = ~(v_w7333_v & v_w7478_v);
	assign v_w6870_v = ~(v_w1821_v & v_w1867_v);
	assign v_o8_v = v_w8037_v ^ v_w8059_v;
	assign v_w7702_v = ~(v_w7700_v | v_w7701_v);
	assign v_w4292_v = ~(v_w4277_v & v_w4280_v);
	assign v_w546_v = v_in32_v ^ v_w545_v;
	assign v_w5172_v = ~(v_w693_v | v_w2194_v);
	assign v_w3484_v = ~(v_w3482_v | v_w3483_v);
	assign v_w3414_v = ~(v_w3412_v | v_w3413_v);
	assign v_w5746_v = ~(v_s272_v & v_w528_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s418_v<=0;
	end
	else
	begin
	v_s418_v<=v_w469_v;
	end
	end
	assign v_w6707_v = ~(v_w6592_v & v_w917_v);
	assign v_w5524_v = ~(v_s189_v & v_w5386_v);
	assign v_w210_v = ~(v_w7874_v & v_w7875_v);
	assign v_w3284_v = ~(v_w3277_v | v_w3283_v);
	assign v_w5678_v = ~(v_s20_v & v_w695_v);
	assign v_w3410_v = ~(v_w3408_v | v_w3409_v);
	assign v_w6728_v = ~(v_w6726_v & v_w6727_v);
	assign v_w1973_v = ~(v_s435_v | v_w1933_v);
	assign v_w3843_v = ~(v_w3839_v & v_w3842_v);
	assign v_w1503_v = ~(v_s300_v ^ v_w1502_v);
	assign v_w2391_v = ~(v_w8220_v);
	assign v_w6137_v = ~(v_w6130_v & v_w6136_v);
	assign v_w5380_v = ~(v_w2916_v | v_w2602_v);
	assign v_w1630_v = ~(v_w1627_v | v_w1629_v);
	assign v_w2167_v = ~(v_w712_v | v_w2166_v);
	assign v_w1524_v = v_w743_v ^ v_w742_v;
	assign v_w2031_v = v_w1100_v ^ v_w2030_v;
	assign v_w7424_v = ~(v_w7419_v & v_w7423_v);
	assign v_w1022_v = ~(v_in23_v & v_w1248_v);
	assign v_w6343_v = ~(v_w6341_v & v_w6342_v);
	assign v_w147_v = v_s138_v & v_w5134_v;
	assign v_w5138_v = ~(v_w5136_v & v_w5137_v);
	assign v_w7288_v = ~(v_w1351_v | v_w680_v);
	assign v_w746_v = ~(v_in16_v ^ v_w1226_v);
	assign v_w5148_v = v_s11_v & v_w5141_v;
	assign v_w1157_v = ~(v_s340_v | v_w1156_v);
	assign v_w2141_v = ~(v_w662_v & v_w1287_v);
	assign v_w118_v = ~(v_w7949_v & v_w7950_v);
	assign v_w2934_v = v_w553_v ^ v_w2933_v;
	assign v_w3489_v = ~(v_w3488_v);
	assign v_w7475_v = ~(v_w7349_v & v_w7474_v);
	assign v_w1893_v = ~(v_w1892_v & v_w917_v);
	assign v_w1582_v = ~(v_w546_v ^ v_w785_v);
	assign v_w3855_v = ~(v_w2406_v & v_w3731_v);
	assign v_w4695_v = ~(v_w674_v & v_s407_v);
	assign v_w7978_v = ~(v_w527_v & v_w7237_v);
	assign v_w5501_v = ~(v_w5499_v | v_w5500_v);
	assign v_w5253_v = ~(v_w2313_v | v_w1_v);
	assign v_w5420_v = ~(v_w5037_v & v_w4825_v);
	assign v_w5251_v = ~(v_w1524_v & v_w5146_v);
	assign v_w3966_v = ~(v_w3774_v & v_w3965_v);
	assign v_w7305_v = ~(v_w7303_v | v_w7304_v);
	assign v_w5227_v = ~(v_s325_v & v_w5141_v);
	assign v_w6225_v = ~(v_w6223_v & v_w6224_v);
	assign v_w6382_v = ~(v_w6379_v ^ v_w6381_v);
	assign v_w7438_v = ~(v_w7434_v & v_w7437_v);
	assign v_w28_v = ~(v_s481_v);
	assign v_w5963_v = ~(v_w5961_v & v_w5962_v);
	assign v_w893_v = ~(v_w1191_v & v_w1278_v);
	assign v_w330_v = ~(v_w5771_v & v_w5782_v);
	assign v_w3088_v = ~(v_w3087_v | v_w557_v);
	assign v_w5681_v = v_w8108_v ^ v_keyinput_32_v;
	assign v_w2931_v = ~(v_w2930_v & v_w569_v);
	assign v_w973_v = ~(v_in22_v ^ v_w1245_v);
	assign v_w3025_v = ~(v_w3012_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s215_v<=0;
	end
	else
	begin
	v_s215_v<=v_w228_v;
	end
	end
	assign v_w5300_v = ~(v_w5124_v & v_w5106_v);
	assign v_w7906_v = ~(v_w651_v & v_w7826_v);
	assign v_w2236_v = ~(v_s170_v | v_w2232_v);
	assign v_w7776_v = ~(v_w7660_v & v_w6787_v);
	assign v_w4454_v = ~(v_w1016_v & v_w2761_v);
	assign v_w1422_v = ~(v_s367_v | v_w1421_v);
	assign v_w462_v = ~(v_w5732_v & v_w5733_v);
	assign v_w7349_v = ~(v_w7344_v & v_w7347_v);
	assign v_w7952_v = ~(v_w527_v & v_w895_v);
	assign v_w4713_v = ~(v_w2342_v | v_w4712_v);
	assign v_w7921_v = ~(v_s274_v & v_w6015_v);
	assign v_w7878_v = ~(v_w651_v & v_w7740_v);
	assign v_w4462_v = ~(v_w4460_v | v_w4461_v);
	assign v_w3711_v = ~(v_w3635_v | v_w3710_v);
	assign v_w5964_v = ~(v_w5959_v | v_w5963_v);
	assign v_w5369_v = ~(v_w683_v & v_w5368_v);
	assign v_w6851_v = ~(v_w1446_v | v_w6571_v);
	assign v_w2027_v = ~(v_w831_v ^ v_w1999_v);
	assign v_w5507_v = ~(v_w683_v & v_w5506_v);
	assign v_w1215_v = ~(v_s93_v & v_w1192_v);
	assign v_w3511_v = ~(v_w2381_v | v_w3510_v);
	assign v_w5425_v = ~(v_w683_v & v_w5424_v);
	assign v_w2554_v = ~(v_w2552_v | v_w2553_v);
	assign v_w5099_v = ~(v_w5098_v & v_w866_v);
	assign v_w1014_v = ~(v_w564_v & v_s76_v);
	assign v_w3048_v = ~(v_w3046_v & v_w3047_v);
	assign v_w124_v = ~(v_w7945_v & v_w7946_v);
	assign v_w1976_v = ~(v_w1975_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s90_v<=0;
	end
	else
	begin
	v_s90_v<=v_w98_v;
	end
	end
	assign v_w8101_v = v_w8100_v ^ v_keyinput_26_v;
	assign v_w3699_v = ~(v_w3518_v | v_w3698_v);
	assign v_w3821_v = ~(v_w3819_v & v_w3820_v);
	assign v_w2168_v = ~(v_w959_v);
	assign v_w2497_v = ~(v_w2495_v & v_w2496_v);
	assign v_w2324_v = ~(v_w8137_v);
	assign v_w7510_v = ~(v_w7508_v & v_w7509_v);
	assign v_w5372_v = ~(v_w5037_v & v_w4944_v);
	assign v_w7212_v = ~(v_w1506_v | v_w7117_v);
	assign v_w4186_v = ~(v_w690_v & v_w4185_v);
	assign v_w3881_v = ~(v_w2588_v | v_w3731_v);
	assign v_w7965_v = ~(v_s27_v & v_w2143_v);
	assign v_w7652_v = v_w529_v & v_w7648_v;
	assign v_w1971_v = ~(v_s475_v & v_w1970_v);
	assign v_w6067_v = ~(v_w6065_v | v_w6066_v);
	assign v_w953_v = ~(v_w951_v & v_w952_v);
	assign v_w2026_v = v_w578_v ^ v_w2015_v;
	assign v_w7841_v = ~(v_s450_v & v_w7667_v);
	assign v_w7879_v = ~(v_s122_v & v_w7876_v);
	assign v_w4129_v = ~(v_w4127_v & v_w4128_v);
	assign v_w4348_v = ~(v_w4347_v & v_w4341_v);
	assign v_w5968_v = ~(v_w5966_v | v_w5967_v);
	assign v_w5866_v = v_w8228_v ^ v_keyinput_112_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s433_v<=0;
	end
	else
	begin
	v_s433_v<=v_w485_v;
	end
	end
	assign v_w6942_v = ~(v_w6938_v | v_w6941_v);
	assign v_w2334_v = ~(v_w568_v | v_w185_v);
	assign v_w605_v = ~(v_w604_v);
	assign v_w7669_v = ~(v_w1835_v & v_w1783_v);
	assign v_w7062_v = ~(v_s273_v & v_w656_v);
	assign v_w8230_v = ~(v_w6029_v | v_w6033_v);
	assign v_w4738_v = ~(v_w4736_v & v_w4737_v);
	assign v_w1444_v = ~(v_w1443_v | v_w808_v);
	assign v_w22_v = ~(v_w5678_v & v_w5679_v);
	assign v_w2656_v = ~(v_w2655_v & v_s384_v);
	assign v_w2072_v = ~(v_w8096_v);
	assign v_w3203_v = ~(v_w2808_v ^ v_w2811_v);
	assign v_w8074_v = v_w1286_v | v_w6608_v;
	assign v_w6970_v = ~(v_w6969_v | v_w6640_v);
	assign v_w3592_v = ~(v_w1007_v | v_w3591_v);
	assign v_w494_v = ~(v_w7827_v & v_w7828_v);
	assign v_w4032_v = ~(v_w688_v | v_w4031_v);
	assign v_w6890_v = ~(v_w1140_v & v_w1459_v);
	assign v_w6532_v = ~(v_w664_v & v_s472_v);
	assign v_w5749_v = ~(v_w662_v & v_w602_v);
	assign v_w1423_v = ~(v_w1422_v | v_w8_v);
	assign v_w3938_v = ~(v_w2753_v | v_w3731_v);
	assign v_o7_v = v_w8039_v ^ v_w8058_v;
	assign v_w1017_v = ~(v_w825_v);
	assign v_w1334_v = ~(v_w1332_v & v_w1333_v);
	assign v_w789_v = ~(v_w989_v);
	assign v_w335_v = ~(v_w5230_v & v_w5231_v);
	assign v_w7108_v = ~(v_w677_v & v_s475_v);
	assign v_w3746_v = ~(v_w3611_v | v_w3731_v);
	assign v_w3170_v = ~(v_w3168_v | v_w3169_v);
	assign v_w1111_v = ~(v_in5_v | v_w1276_v);
	assign v_w3174_v = ~(v_w3171_v | v_w3173_v);
	assign v_w798_v = ~(v_w1725_v | v_w998_v);
	assign v_w5314_v = ~(v_s240_v & v_w5293_v);
	assign v_w5636_v = ~(v_s213_v & v_w695_v);
	assign v_w4892_v = ~(v_w2448_v & v_w2937_v);
	assign v_w8046_v = ~(v_w7984_v | v_w8045_v);
	assign v_w4782_v = ~(v_w4781_v | v_w4589_v);
	assign v_w4278_v = ~(v_w2930_v & v_s350_v);
	assign v_w1035_v = ~(v_w531_v & v_s250_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s410_v<=0;
	end
	else
	begin
	v_s410_v<=v_w459_v;
	end
	end
	assign v_w5326_v = ~(v_w5324_v | v_w5325_v);
	assign v_w4939_v = ~(v_w2347_v & v_w2840_v);
	assign v_w3159_v = ~(v_w2840_v & v_w2634_v);
	assign v_w5960_v = ~(v_w986_v ^ v_w2023_v);
	assign v_w471_v = ~(v_w7850_v & v_w7851_v);
	assign v_w863_v = ~(v_w2294_v | v_w1703_v);
	assign v_w3460_v = v_w8167_v ^ v_keyinput_72_v;
	assign v_w5858_v = ~(v_w600_v & v_w2063_v);
	assign v_w1327_v = ~(v_w1067_v & v_w1323_v);
	assign v_w2469_v = ~(v_w2459_v | v_w2468_v);
	assign v_w165_v = ~(v_w3335_v & v_w3337_v);
	assign v_w295_v = ~(v_s495_v);
	assign v_w8068_v = v_w8067_v ^ v_keyinput_3_v;
	assign v_w1433_v = ~(v_w1429_v | v_w1432_v);
	assign v_w4028_v = v_w8175_v ^ v_keyinput_79_v;
	assign v_w955_v = ~(v_w844_v | v_w954_v);
	assign v_w8124_v = ~(v_w3960_v | v_w3963_v);
	assign v_w8130_v = v_w2635_v | v_w2581_v;
	assign v_w5618_v = ~(v_s5_v & v_w676_v);
	assign v_w7630_v = ~(v_w7595_v & v_w7629_v);
	assign v_w2319_v = ~(v_w2293_v | v_w1561_v);
	assign v_w4859_v = ~(v_w2952_v & v_w2347_v);
	assign v_w2444_v = ~(v_w2392_v | v_w2443_v);
	assign v_w1421_v = ~(v_w720_v | v_w8_v);
	assign v_w8025_v = ~(v_s461_v ^ v_s311_v);
	assign v_w7139_v = ~(v_w7118_v & v_w1299_v);
	assign v_w2376_v = ~(v_w2358_v & v_s294_v);
	assign v_w3842_v = ~(v_w3840_v & v_w3841_v);
	assign v_w1080_v = ~(v_w3200_v | v_w3201_v);
	assign v_w4655_v = ~(v_w2690_v & v_w2369_v);
	assign v_w6929_v = ~(v_w1642_v | v_w1797_v);
	assign v_w6016_v = ~(v_w890_v | v_w6015_v);
	assign v_w833_v = ~(v_w1517_v | v_w808_v);
	assign v_w1216_v = ~(v_w612_v & v_s95_v);
	assign v_w6401_v = ~(v_w6398_v ^ v_w6400_v);
	assign v_w63_v = v_s55_v & v_w7107_v;
	assign v_w4702_v = ~(v_w2448_v & v_w2722_v);
	assign v_w5413_v = ~(v_w5411_v | v_w5412_v);
	assign v_w2596_v = ~(v_w2569_v ^ v_w2595_v);
	assign v_w1623_v = ~(v_w1621_v & v_w1622_v);
	assign v_w1957_v = ~(v_s74_v | v_s73_v);
	assign v_w6857_v = ~(v_w1680_v);
	assign v_w1521_v = v_s287_v ^ v_w1148_v;
	assign v_w7150_v = ~(v_w7118_v & v_w1339_v);
	assign v_w3917_v = ~(v_w3916_v & v_w956_v);
	assign v_w5512_v = ~(v_w4863_v | v_w4622_v);
	assign v_w774_v = ~(v_w772_v | v_w773_v);
	assign v_w3840_v = ~(v_w3735_v & v_w2367_v);
	assign v_w2348_v = ~(v_w2346_v & v_w2347_v);
	assign v_w742_v = v_in29_v ^ v_w1268_v;
	assign v_w8168_v = v_w8035_v ^ v_w8060_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s323_v<=0;
	end
	else
	begin
	v_s323_v<=v_w349_v;
	end
	end
	assign v_w1249_v = v_in23_v ^ v_w1248_v;
	assign v_w3179_v = ~(v_w3031_v & v_w2634_v);
	assign v_w5174_v = ~(v_w8170_v);
	assign v_w1604_v = ~(v_w1601_v | v_w1603_v);
	assign v_w4058_v = ~(v_s260_v & v_w693_v);
	assign v_w4422_v = ~(v_w1069_v & v_w4421_v);
	assign v_w7434_v = ~(v_w7379_v & v_w7433_v);
	assign v_w2971_v = ~(v_w582_v | v_w583_v);
	assign v_w6508_v = ~(v_s102_v & v_w888_v);
	assign v_w2912_v = ~(v_w2902_v & v_w2911_v);
	assign v_w5383_v = ~(v_w5382_v | v_w4929_v);
	assign v_w503_v = ~(v_w7840_v & v_w7841_v);
	assign v_w5509_v = ~(v_w4625_v & v_w5126_v);
	assign v_w134_v = ~(v_w5194_v & v_w5195_v);
	assign v_w7464_v = ~(v_w7456_v & v_w7463_v);
	assign v_w5329_v = ~(v_s230_v & v_w5293_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s221_v<=0;
	end
	else
	begin
	v_s221_v<=v_w234_v;
	end
	end
	assign v_w8107_v = v_w8106_v ^ v_keyinput_31_v;
	assign v_w3516_v = ~(v_w3515_v);
	assign v_w5076_v = ~(v_w2400_v | v_w2370_v);
	assign v_w1373_v = ~(v_w1369_v | v_w1372_v);
	assign v_w5339_v = ~(v_w2601_v & v_w2558_v);
	assign v_w2502_v = ~(v_w2331_v | v_w617_v);
	assign v_w691_v = ~(v_w2266_v & v_w1037_v);
	assign v_w5775_v = ~(v_w2031_v & v_w728_v);
	assign v_w2079_v = ~(v_w1350_v | v_w2078_v);
	assign v_w3808_v = v_w3804_v | v_w3807_v;
	assign v_w7046_v = ~(v_w7045_v & v_w1915_v);
	assign v_w7042_v = ~(v_w7038_v | v_w7041_v);
	assign v_w6313_v = ~(v_w6301_v | v_w6312_v);
	assign v_w5453_v = ~(v_w2601_v & v_w760_v);
	assign v_w3107_v = ~(v_w3084_v ^ v_w3106_v);
	assign v_w2873_v = ~(v_w2871_v & v_w2872_v);
	assign v_w6306_v = ~(v_w6304_v ^ v_w6305_v);
	assign v_w3896_v = ~(v_w3822_v & v_w3895_v);
	assign v_w6222_v = ~(v_w6208_v | v_w6221_v);
	assign v_w6517_v = ~(v_w6516_v | v_w6015_v);
	assign v_w1425_v = ~(v_w1424_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s485_v<=0;
	end
	else
	begin
	v_s485_v<=v_w47_v;
	end
	end
	assign v_w1094_v = ~(v_w1092_v | v_w1093_v);
	assign v_w6817_v = ~(v_w6807_v | v_w6816_v);
	assign v_w167_v = ~(v_w5908_v & v_w5909_v);
	assign v_w7455_v = ~(v_w7439_v & v_w7454_v);
	assign v_w6907_v = ~(v_w1140_v & v_w1638_v);
	assign v_w4640_v = ~(v_w2265_v & v_w755_v);
	assign v_w1547_v = ~(v_s272_v | v_w1180_v);
	assign v_w1311_v = ~(v_w1309_v);
	assign v_w1363_v = ~(v_w1362_v);
	assign v_w6721_v = ~(v_w6719_v | v_w6720_v);
	assign v_w3977_v = ~(v_w3975_v & v_w3976_v);
	assign v_w2446_v = ~(v_w2445_v & v_w878_v);
	assign v_w4903_v = v_w572_v ^ v_w4404_v;
	assign v_w1068_v = ~(v_w3486_v & v_w3487_v);
	assign v_w6824_v = ~(v_w1417_v | v_w1419_v);
	assign v_w1539_v = ~(v_s269_v ^ v_w1538_v);
	assign v_w5486_v = ~(v_w5483_v & v_w5485_v);
	assign v_w8067_v = v_w2471_v ^ v_w2441_v;
	assign v_w2799_v = ~(v_w2797_v | v_w2798_v);
	assign v_w7626_v = ~(v_w1286_v | v_w1003_v);
	assign v_w7420_v = v_w5905_v ^ v_w1781_v;
	assign v_w252_v = ~(v_w5564_v & v_w5565_v);
	assign v_w592_v = ~(v_w2354_v);
	assign v_w360_v = ~(v_w4246_v & v_w4256_v);
	assign v_w7736_v = ~(v_s196_v & v_w7667_v);
	assign v_w3669_v = ~(v_w3636_v & v_w3668_v);
	assign v_w501_v = ~(v_w2114_v & v_w869_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s482_v<=0;
	end
	else
	begin
	v_s482_v<=v_w33_v;
	end
	end
	assign v_w7158_v = ~(v_w7118_v & v_w1715_v);
	assign v_w46_v = ~(v_w5606_v & v_w5607_v);
	assign v_w5282_v = ~(v_w5281_v ^ v_w3678_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s235_v<=0;
	end
	else
	begin
	v_s235_v<=v_w248_v;
	end
	end
	assign v_w6471_v = ~(v_w6469_v & v_w6470_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s26_v<=0;
	end
	else
	begin
	v_s26_v<=v_w29_v;
	end
	end
	assign v_w4534_v = v_w3556_v & v_w3552_v;
	assign v_w5765_v = ~(v_w5761_v | v_w5764_v);
	assign v_w4509_v = ~(v_w4449_v & v_w4508_v);
	assign v_w7831_v = ~(v_w7830_v | v_w6632_v);
	assign v_w2151_v = ~(v_s276_v | v_s275_v);
	assign v_w6085_v = ~(v_w1579_v | v_w6062_v);
	assign v_w8140_v = ~(v_w4448_v & v_w4513_v);
	assign v_w2278_v = ~(v_w947_v & v_w2153_v);
	assign v_w7444_v = ~(v_w1856_v | v_w680_v);
	assign v_w4491_v = ~(v_w4489_v | v_w4490_v);
	assign v_w3725_v = ~(v_w3724_v & v_w3489_v);
	assign v_w1393_v = ~(v_w613_v & v_w1392_v);
	assign v_w6077_v = v_s246_v ^ v_w1557_v;
	assign v_w1597_v = ~(v_w1596_v & v_w980_v);
	assign v_w5903_v = ~(v_w2137_v & v_w1834_v);
	assign v_w1406_v = ~(v_s373_v & v_w562_v);
	assign v_w4520_v = ~(v_w4518_v | v_w4519_v);
	assign v_w1845_v = ~(v_w950_v & v_w1028_v);
	assign v_w584_v = ~(v_w582_v ^ v_w583_v);
	assign v_w4428_v = ~(v_w4426_v | v_w4427_v);
	assign v_w1622_v = ~(v_w666_v & v_s204_v);
	assign v_w3150_v = ~(v_w3149_v & v_w3126_v);
	assign v_w7696_v = ~(v_w8118_v);
	assign v_w5597_v = ~(v_w5555_v & v_w5460_v);
	assign v_w1149_v = v_s287_v | v_w1148_v;
	assign v_w5428_v = ~(v_w5037_v & v_w4796_v);
	assign v_w3992_v = ~(v_w3984_v | v_w3991_v);
	assign v_w2721_v = ~(v_w2355_v & v_s83_v);
	assign v_w1370_v = ~(v_w1052_v & v_s98_v);
	assign v_w497_v = ~(v_s518_v);
	assign v_w1817_v = ~(v_w847_v);
	assign v_w3697_v = ~(v_w3695_v | v_w3696_v);
	assign v_w6886_v = ~(v_w1094_v | v_w6579_v);
	assign v_w7025_v = ~(v_w1521_v | v_w6571_v);
	assign v_w4612_v = ~(v_w4526_v | v_w4604_v);
	assign v_w7181_v = ~(v_w7179_v | v_w7180_v);
	assign v_w8109_v = v_w6419_v & v_w6423_v;
	assign v_w4232_v = ~(v_w690_v & v_w4231_v);
	assign v_w6050_v = ~(v_w6047_v | v_w6049_v);
	assign v_w7246_v = ~(v_w687_v & v_w7245_v);
	assign v_w2466_v = ~(v_w2460_v | v_w2465_v);
	assign v_w4791_v = ~(v_w4785_v & v_w4790_v);
	assign v_w1603_v = ~(v_w1602_v | v_w1180_v);
	assign v_w567_v = ~(v_w566_v);
	assign v_w5538_v = ~(v_w1069_v | v_w2602_v);
	assign v_w3497_v = ~(v_w3496_v & v_w2431_v);
	assign v_w490_v = ~(v_w5821_v & v_w5827_v);
	assign v_w2589_v = ~(v_w2588_v | v_w557_v);
	assign v_w6336_v = ~(v_w5948_v & v_w6335_v);
	assign v_w3246_v = ~(v_w3245_v & v_w2944_v);
	assign v_w7284_v = ~(v_w1363_v | v_w680_v);
	assign v_w1875_v = ~(v_w1436_v & v_w1091_v);
	assign v_w2212_v = ~(v_w2210_v & v_w2211_v);
	assign v_w5839_v = ~(v_w5837_v | v_w5838_v);
	assign v_w2252_v = ~(v_w2248_v & v_w2251_v);
	assign v_w7186_v = ~(v_s120_v & v_w7112_v);
	assign v_w320_v = ~(v_w5632_v & v_w5633_v);
	assign v_w7957_v = ~(v_s82_v & v_w2143_v);
	assign v_w2401_v = ~(v_w2400_v | v_w2317_v);
	assign v_w2699_v = ~(v_w699_v & v_s422_v);
	assign v_w2571_v = v_s310_v ^ v_w2551_v;
	assign v_w2824_v = ~(v_w2823_v & v_w569_v);
	assign v_w6827_v = ~(v_w6823_v & v_w6826_v);
	assign v_w1400_v = ~(v_w875_v & v_s355_v);
	assign v_w2270_v = ~(v_w2267_v | v_w2269_v);
	assign v_w3124_v = ~(v_w584_v ^ v_w2969_v);
	assign v_w6876_v = ~(v_w8250_v);
	assign v_w6993_v = ~(v_w1496_v | v_w6571_v);
	assign v_w540_v = ~(v_in29_v & v_w1268_v);
	assign v_w2593_v = v_w552_v ^ v_w2592_v;
	assign v_w6360_v = ~(v_w6358_v & v_w6359_v);
	assign v_w640_v = ~(v_w2913_v & v_w2918_v);
	assign v_w6542_v = v_s402_v ^ v_w1772_v;
	assign v_w3600_v = ~(v_w3586_v & v_w3599_v);
	assign v_w3439_v = ~(v_w2773_v | v_w2620_v);
	assign v_w2452_v = ~(v_w674_v | v_w2451_v);
	assign v_w6014_v = ~(v_w659_v & v_w396_v);
	assign v_w4741_v = ~(v_w4502_v ^ v_w3633_v);
	assign v_w7639_v = ~(v_w7635_v & v_w7638_v);
	assign v_w3228_v = ~(v_w3226_v & v_w3227_v);
	assign v_w7566_v = ~(v_w5905_v | v_w7565_v);
	assign v_w4160_v = v_s229_v ^ v_w4153_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s299_v<=0;
	end
	else
	begin
	v_s299_v<=v_w321_v;
	end
	end
	assign v_w2832_v = ~(v_w558_v & v_w2831_v);
	assign v_w3858_v = ~(v_w2327_v & v_w881_v);
	assign v_w1986_v = ~(v_w1782_v | v_w883_v);
	assign v_w5566_v = ~(v_s231_v & v_w676_v);
	assign v_w7757_v = ~(v_w7756_v | v_w6845_v);
	assign v_w7296_v = ~(v_w687_v | v_w1725_v);
	assign v_w8020_v = ~(v_w8018_v | v_w8019_v);
	assign v_w5569_v = ~(v_w675_v & v_w5345_v);
	assign v_w433_v = ~(v_w3257_v & v_w3263_v);
	assign v_w7354_v = ~(v_w687_v | v_w1126_v);
	assign v_w3352_v = ~(v_s360_v & v_w693_v);
	assign v_w3223_v = ~(v_s260_v & v_w3222_v);
	assign v_w3121_v = ~(v_w2639_v);
	assign v_w1316_v = v_s436_v ^ v_w1167_v;
	assign v_w6256_v = v_w6251_v ^ v_w6255_v;
	assign v_w2183_v = ~(v_w2181_v | v_w2182_v);
	assign v_w2927_v = ~(v_w2926_v | v_w557_v);
	assign v_w627_v = ~(v_w2058_v & v_w1435_v);
	assign v_w444_v = ~(v_w4386_v & v_w4396_v);
	assign v_w4268_v = ~(v_w2929_v ^ v_s352_v);
	assign v_w1011_v = ~(v_w1009_v | v_w1010_v);
	assign v_w5994_v = ~(v_w2113_v & v_w5993_v);
	assign v_w1690_v = ~(v_w1404_v | v_w1689_v);
	assign v_w5296_v = ~(v_w5131_v & v_w5295_v);
	assign v_w595_v = ~(v_w1561_v | v_w808_v);
	assign v_w95_v = ~(v_w7917_v & v_w7918_v);
	assign v_w1049_v = v_in14_v ^ v_w1220_v;
	assign v_w2271_v = ~(v_w2270_v & v_w2152_v);
	assign v_w7345_v = ~(v_w687_v | v_w1094_v);
	assign v_w7559_v = ~(v_w8087_v);
	assign v_w4293_v = ~(v_w4291_v & v_w4292_v);
	assign v_w73_v = v_s65_v & v_w7107_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s152_v<=0;
	end
	else
	begin
	v_s152_v<=v_w161_v;
	end
	end
	assign v_w2615_v = ~(v_w2361_v | v_w2614_v);
	assign v_w4836_v = ~(v_w4826_v & v_w4835_v);
	assign v_w4776_v = ~(v_w3338_v & v_w2369_v);
	assign v_w2015_v = ~(v_w567_v ^ v_w1999_v);
	assign v_w1530_v = ~(v_w875_v & v_s286_v);
	assign v_w2765_v = ~(v_w2760_v | v_w2764_v);
	assign v_w8004_v = v_s280_v ^ v_s457_v;
	assign v_w5388_v = ~(v_w4906_v & v_w5126_v);
	assign v_w5633_v = ~(v_w420_v & v_w2367_v);
	assign v_w7826_v = ~(v_w7824_v & v_w7825_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s88_v<=0;
	end
	else
	begin
	v_s88_v<=v_w96_v;
	end
	end
	assign v_w6719_v = ~(v_w6717_v & v_w6718_v);
	assign v_w6356_v = ~(v_w6352_v ^ v_w6355_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s55_v<=0;
	end
	else
	begin
	v_s55_v<=v_w63_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s137_v<=0;
	end
	else
	begin
	v_s137_v<=v_w146_v;
	end
	end
	assign v_w3153_v = ~(v_w3109_v & v_w2910_v);
	assign v_w7223_v = ~(v_w1539_v | v_w528_v);
	assign v_w6234_v = ~(v_w5772_v & v_w6233_v);
	assign v_w2586_v = ~(v_w2484_v & v_w2585_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s432_v<=0;
	end
	else
	begin
	v_s432_v<=v_w483_v;
	end
	end
	assign v_w7361_v = ~(v_w687_v | v_w1656_v);
	assign v_w2646_v = ~(v_w2645_v & v_s360_v);
	assign v_w4207_v = ~(v_w2822_v ^ v_s316_v);
	assign v_w1904_v = ~(v_w1901_v & v_w1903_v);
	assign v_w2383_v = ~(v_w2382_v);
	assign v_w748_v = ~(v_w746_v | v_w747_v);
	assign v_w50_v = ~(v_w5602_v & v_w5603_v);
	assign v_w2137_v = ~(v_w661_v | v_w2136_v);
	assign v_w1808_v = ~(v_w1309_v | v_w1064_v);
	assign v_w4873_v = ~(v_w4867_v | v_w4589_v);
	assign v_w3510_v = ~(v_w3509_v);
	assign v_w3672_v = ~(v_w781_v | v_w3671_v);
	assign v_w5572_v = ~(v_s212_v & v_w676_v);
	assign v_w3341_v = ~(v_w3339_v & v_w3340_v);
	assign v_w5068_v = ~(v_w5066_v & v_w5067_v);
	assign v_w1874_v = ~(v_w1872_v & v_w1873_v);
	assign v_w8249_v = v_w6873_v & v_w6875_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s163_v<=0;
	end
	else
	begin
	v_s163_v<=v_w172_v;
	end
	end
	assign v_w1671_v = ~(v_w666_v & v_s121_v);
	assign v_w3061_v = ~(v_w558_v & v_w3060_v);
	assign v_w1161_v = v_s343_v | v_w1160_v;
	assign v_w1516_v = ~(v_w562_v & v_s232_v);
	assign v_w5087_v = ~(v_w5084_v | v_w5086_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s92_v<=0;
	end
	else
	begin
	v_s92_v<=v_w100_v;
	end
	end
	assign v_w7830_v = ~(v_w7829_v | v_w1919_v);
	assign v_w8162_v = ~(v_w6388_v & v_w659_v);
	assign v_w6599_v = ~(v_w2102_v ^ v_w6598_v);
	assign v_w7790_v = ~(v_w654_v & v_w7789_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s136_v<=0;
	end
	else
	begin
	v_s136_v<=v_w145_v;
	end
	end
	assign v_w6838_v = ~(v_w6837_v & v_w1915_v);
	assign v_w7190_v = ~(v_s193_v & v_w7112_v);
	assign v_w5979_v = ~(v_w5977_v & v_w5978_v);
	assign v_w171_v = ~(v_w5210_v & v_w5211_v);
	assign v_w810_v = ~(v_w2713_v | v_w764_v);
	assign v_w6727_v = v_w6571_v | v_w1355_v;
	assign v_w4935_v = ~(v_w4932_v | v_w4934_v);
	assign v_w2224_v = ~(v_s133_v | v_s132_v);
	assign v_w8158_v = ~(v_w1614_v & v_w1615_v);
	assign v_w7269_v = ~(v_w687_v & v_w1065_v);
	assign v_w4010_v = ~(v_w3741_v & v_w4009_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s291_v<=0;
	end
	else
	begin
	v_s291_v<=v_w311_v;
	end
	end
	assign v_w6066_v = ~(v_w6018_v | v_w1579_v);
	assign v_w3035_v = ~(v_w3030_v | v_w3034_v);
	assign v_w6006_v = ~(v_w6005_v & v_w2113_v);
	assign v_w2899_v = ~(v_w2895_v | v_w2898_v);
	assign v_w2264_v = ~(v_w2263_v & v_w673_v);
	assign v_w8040_v = ~(v_w7990_v | v_w8039_v);
	assign v_w7981_v = ~(v_s471_v | v_s390_v);
	assign v_w683_v = v_w681_v & v_w682_v;
	assign v_w2481_v = ~(v_w2479_v & v_w2480_v);
	assign v_w6759_v = ~(v_w6757_v & v_w6758_v);
	assign v_w1469_v = ~(v_w1466_v | v_w1468_v);
	assign v_w2234_v = ~(v_w865_v & v_w555_v);
	assign v_w2964_v = ~(v_w2957_v | v_w2963_v);
	assign v_w4034_v = ~(v_w4032_v | v_w4033_v);
	assign v_w4937_v = ~(v_w2856_v | v_w2264_v);
	assign v_w3139_v = ~(v_w3109_v & v_w2706_v);
	assign v_w256_v = ~(v_w7685_v & v_w7686_v);
	assign v_w3461_v = ~(v_w855_v & v_w3460_v);
	assign v_w1929_v = ~(v_w1928_v ^ v_s12_v);
	assign v_w126_v = ~(v_w5586_v & v_w5587_v);
	assign v_w5091_v = ~(v_w5089_v & v_w5090_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s464_v<=0;
	end
	else
	begin
	v_s464_v<=v_w517_v;
	end
	end
	assign v_w3825_v = ~(v_w3823_v | v_w3824_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s197_v<=0;
	end
	else
	begin
	v_s197_v<=v_w210_v;
	end
	end
	assign v_w3744_v = ~(v_w881_v | v_w963_v);
	assign v_w414_v = ~(v_w4824_v & v_w4837_v);
	assign v_w6505_v = ~(v_w6503_v | v_w6504_v);
	assign v_w4066_v = ~(v_w4059_v | v_w4065_v);
	assign v_w3144_v = ~(v_w3141_v | v_w3143_v);
	assign v_w3827_v = ~(v_w3521_v | v_w3731_v);
	assign v_w7653_v = ~(v_s433_v & v_w1971_v);
	assign v_w2941_v = v_w2888_v & v_w2892_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s510_v<=0;
	end
	else
	begin
	v_s510_v<=v_w400_v;
	end
	end
	assign v_w3218_v = ~(v_w3109_v & v_w1131_v);
	assign v_w6333_v = ~(v_s338_v ^ v_w6332_v);
	assign v_w6054_v = ~(v_w6042_v | v_w1579_v);
	assign v_w7017_v = ~(v_w7016_v | v_w6594_v);
	assign v_o5_v = v_w8043_v ^ v_w8056_v;
	assign v_w79_v = v_s71_v & v_w7107_v;
	assign v_w2810_v = ~(v_w2484_v & v_w2618_v);
	assign v_w1855_v = ~(v_w923_v & v_w1854_v);
	assign v_w7994_v = v_s465_v & v_s332_v;
	assign v_w7497_v = ~(v_w7309_v & v_w7496_v);
	assign v_w6687_v = ~(v_w6685_v & v_w6686_v);
	assign v_w2512_v = ~(v_w2406_v | v_w557_v);
	assign v_w2173_v = ~(v_w2169_v | v_w2172_v);
	assign v_w2622_v = ~(v_w2609_v | v_w2621_v);
	assign v_w2374_v = ~(v_w2372_v & v_w2373_v);
	assign v_w2869_v = ~(v_w2867_v & v_w2868_v);
	assign v_w6656_v = ~(v_w6654_v & v_w6655_v);
	assign v_w1568_v = v_w1051_v & v_s357_v;
	assign v_w4720_v = ~(v_w4718_v & v_w4719_v);
	assign v_w4908_v = v_w4549_v ^ v_w3641_v;
	assign v_w6746_v = ~(v_w884_v & v_w6745_v);
	assign v_w2443_v = ~(v_w2438_v | v_w2442_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s516_v<=0;
	end
	else
	begin
	v_s516_v<=v_w460_v;
	end
	end
	assign v_w692_v = ~(v_w691_v | v_w689_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s227_v<=0;
	end
	else
	begin
	v_s227_v<=v_w240_v;
	end
	end
	assign v_w4857_v = ~(v_w4854_v | v_w4856_v);
	assign v_w4715_v = v_w2261_v | v_w2718_v;
	assign v_w729_v = ~(v_w1551_v | v_w1554_v);
	assign v_w2419_v = ~(v_w2335_v);
	assign v_w4896_v = ~(v_w4889_v & v_w4895_v);
	assign v_w3039_v = ~(v_w1078_v | v_w616_v);
	assign v_w6659_v = ~(v_w1809_v | v_w1808_v);
	assign v_w1351_v = ~(v_w1350_v);
	assign v_w2428_v = ~(v_w2427_v);
	assign v_w3476_v = ~(v_w3474_v | v_w3475_v);
	assign v_w6973_v = ~(v_w6592_v & v_w919_v);
	assign v_w5232_v = ~(v_w1476_v | v_w5145_v);
	assign v_w2249_v = ~(v_w2164_v | v_w2191_v);
	assign v_w476_v = ~(v_w4428_v & v_w4432_v);
	assign v_w8049_v = ~(v_w7981_v | v_w8048_v);
	assign v_w6553_v = ~(v_s102_v & v_w1701_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s340_v<=0;
	end
	else
	begin
	v_s340_v<=v_w371_v;
	end
	end
	assign v_w4092_v = ~(v_w4090_v & v_w4091_v);
	assign v_w6552_v = ~(v_w6029_v | v_w6551_v);
	assign v_w2515_v = v_w2514_v ^ v_w552_v;
	assign v_w3328_v = ~(v_w3324_v | v_w3327_v);
	assign v_w2152_v = ~(v_w2150_v & v_w2151_v);
	assign v_w5316_v = ~(v_w5056_v & v_w5126_v);
	assign v_w7508_v = ~(v_w7506_v | v_w7507_v);
	assign v_w1758_v = ~(v_w870_v & v_w1757_v);
	assign v_w1476_v = v_w977_v ^ v_w976_v;
	assign v_w4796_v = v_w4409_v ^ v_w1011_v;
	assign v_w5244_v = ~(v_w693_v | v_w2289_v);
	assign v_w1921_v = ~(v_w1917_v | v_w1920_v);
	assign v_w3740_v = ~(v_w3738_v | v_w3739_v);
	assign v_w7421_v = ~(v_w7420_v & v_w686_v);
	assign v_w4964_v = ~(v_w4961_v | v_w4963_v);
	assign v_w7166_v = ~(v_s393_v & v_w7113_v);
	assign v_w3479_v = ~(v_s8_v & v_w564_v);
	assign v_w6924_v = ~(v_w1624_v | v_w6608_v);
	assign v_w3748_v = ~(v_w3746_v | v_w3747_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s288_v<=0;
	end
	else
	begin
	v_s288_v<=v_w308_v;
	end
	end
	assign v_w6745_v = ~(v_w6744_v);
	assign v_w4571_v = ~(v_w4533_v | v_w4570_v);
	assign v_w2425_v = ~(v_w2423_v & v_w2424_v);
	assign v_w6893_v = ~(v_w6891_v | v_w6892_v);
	assign v_w4456_v = v_w3490_v & v_w3553_v;
	assign v_w3135_v = ~(v_w3133_v | v_w3134_v);
	assign v_w4029_v = ~(v_w3623_v | v_w4028_v);
	assign v_w4530_v = ~(v_w4446_v | v_w4529_v);
	assign v_w371_v = ~(v_w5926_v & v_w5933_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s169_v<=0;
	end
	else
	begin
	v_s169_v<=v_w179_v;
	end
	end
	assign v_w1698_v = ~(v_w1695_v & v_w1697_v);
	assign v_w5191_v = ~(v_s99_v & v_w5141_v);
	assign v_w4706_v = ~(v_w4705_v | v_w4589_v);
	assign v_w1434_v = ~(v_w1052_v & v_s114_v);
	assign v_w7182_v = ~(v_s366_v & v_w7112_v);
	assign v_w3689_v = ~(v_w3688_v & v_w3482_v);
	assign v_w565_v = v_w563_v;
	assign v_w533_v = ~(v_s521_v);
	assign v_w5949_v = ~(v_w5947_v & v_w5948_v);
	assign v_w4440_v = ~(v_w3114_v & v_w2347_v);
	assign v_w4662_v = ~(v_w4659_v | v_w4661_v);
	assign v_w6735_v = ~(v_w6734_v ^ v_w1887_v);
	assign v_w2797_v = ~(v_s217_v | v_w2796_v);
	assign v_w1887_v = ~(v_w1364_v & v_w1730_v);
	assign v_w2186_v = v_w712_v & v_w2154_v;
	assign v_w5510_v = ~(v_w2601_v & v_w871_v);
	assign v_w1735_v = ~(v_w1734_v & v_w1350_v);
	assign v_w7679_v = ~(v_w654_v & v_w7678_v);
	assign v_w448_v = ~(v_w5974_v & v_w5976_v);
	assign v_w3175_v = ~(v_s380_v & v_w1_v);
	assign v_w6842_v = v_w1687_v ^ v_w1873_v;
	assign v_w7582_v = ~(v_w1736_v | v_w7581_v);
	assign v_w2774_v = ~(v_w2773_v | v_w538_v);
	assign v_w3448_v = ~(v_s192_v & v_w699_v);
	assign v_w4202_v = ~(v_w4200_v & v_w4201_v);
	assign v_w3536_v = ~(v_w3535_v);
	assign v_w4778_v = ~(v_w4777_v & v_w878_v);
	assign v_w7815_v = ~(v_w654_v & v_w7814_v);
	assign v_w2143_v = ~(v_w2118_v & v_w1969_v);
	assign v_w5856_v = ~(v_w5854_v | v_w5855_v);
	assign v_w7634_v = ~(v_w7631_v | v_w7633_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s9_v<=0;
	end
	else
	begin
	v_s9_v<=v_w10_v;
	end
	end
	assign v_w7837_v = ~(v_w1803_v | v_w1782_v);
	assign v_w1288_v = v_w805_v ^ v_w1060_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s129_v<=0;
	end
	else
	begin
	v_s129_v<=v_w138_v;
	end
	end
	assign v_w959_v = ~(v_s162_v | v_w927_v);
	assign v_w1102_v = ~(v_in30_v & v_w1271_v);
	assign v_w7726_v = ~(v_w6934_v | v_w7725_v);
	assign v_w8203_v = v_w8202_v ^ v_keyinput_97_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s51_v<=0;
	end
	else
	begin
	v_s51_v<=v_w59_v;
	end
	end
	assign v_w6445_v = v_w1424_v ^ v_w6444_v;
	assign v_w5459_v = ~(v_w5457_v | v_w5458_v);
	assign v_w4910_v = ~(v_w2447_v & v_w2910_v);
	assign v_w5288_v = ~(v_w5278_v | v_w5287_v);
	assign v_w1407_v = v_s374_v ^ v_w1388_v;
	assign v_w5097_v = v_w2419_v ^ v_w2331_v;
	assign v_w4264_v = ~(v_w4263_v & v_w690_v);
	assign v_w6462_v = ~(v_w657_v & v_s406_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s412_v<=0;
	end
	else
	begin
	v_s412_v<=v_w463_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s324_v<=0;
	end
	else
	begin
	v_s324_v<=v_w350_v;
	end
	end
	assign v_w7643_v = ~(v_w7593_v | v_w7642_v);
	assign v_w5271_v = v_w4421_v ^ v_w1069_v;
	assign v_w8234_v = v_w8233_v ^ v_keyinput_116_v;
	assign v_w3379_v = ~(v_s328_v & v_w693_v);
	assign v_w513_v = ~(v_w6194_v & v_w6206_v);
	assign v_w3939_v = ~(v_w3937_v | v_w3938_v);
	assign v_w5312_v = ~(v_w5087_v & v_w5311_v);
	assign v_w7239_v = v_w7238_v ^ v_keyinput_65_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s477_v<=0;
	end
	else
	begin
	v_s477_v<=v_w532_v;
	end
	end
	assign v_w8094_v = ~(v_w3763_v & v_w3766_v);
	assign v_w2513_v = ~(v_w2326_v | v_w617_v);
	assign v_w4215_v = ~(v_w4191_v | v_w4189_v);
	assign v_w2695_v = ~(v_w2484_v & v_w2690_v);
	assign v_w1143_v = ~(v_w1192_v | v_w3464_v);
	assign v_w2545_v = ~(v_w2541_v | v_w2544_v);
	assign v_w3469_v = ~(v_w3468_v);
	assign v_w1198_v = ~(v_w1196_v & v_w1197_v);
	assign v_w2740_v = ~(v_w2730_v & v_w2739_v);
	assign v_w3962_v = ~(v_w3567_v | v_w3735_v);
	assign v_w1356_v = ~(v_w1355_v | v_w1180_v);
	assign v_w2782_v = ~(v_w2781_v & v_w844_v);
	assign v_w2060_v = ~(v_w1021_v ^ v_w1999_v);
	assign v_w4600_v = ~(v_w2342_v | v_w4599_v);
	assign v_w7968_v = ~(v_w527_v & v_w1297_v);
	assign v_w3090_v = ~(v_w2358_v & v_s428_v);
	assign v_w5809_v = ~(v_w5807_v & v_w5808_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s283_v<=0;
	end
	else
	begin
	v_s283_v<=v_w302_v;
	end
	end
	assign v_w6895_v = ~(v_w6894_v | v_w6594_v);
	assign v_w5956_v = ~(v_w5955_v & v_w5703_v);
	assign v_w6803_v = v_w1689_v ^ v_w6802_v;
	assign v_w7183_v = ~(v_w1667_v | v_w529_v);
	assign v_w4226_v = ~(v_w2851_v ^ v_s329_v);
	assign v_w5936_v = ~(v_w662_v & v_w1362_v);
	assign v_w3989_v = ~(v_w3587_v & v_w881_v);
	assign v_w3612_v = ~(v_w3611_v | v_w963_v);
	assign v_w8163_v = ~(v_w6988_v & v_w655_v);
	assign v_w7852_v = ~(v_s357_v & v_w1993_v);
	assign v_w2075_v = ~(v_w2073_v | v_w2074_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s382_v<=0;
	end
	else
	begin
	v_s382_v<=v_w428_v;
	end
	end
	assign v_w3155_v = ~(v_w3151_v | v_w3154_v);
	assign v_w8021_v = ~(v_w8001_v | v_w8020_v);
	assign v_w290_v = ~(v_w5752_v & v_w5756_v);
	assign v_w6537_v = ~(v_w1700_v | v_w6029_v);
	assign v_w3583_v = ~(v_w3582_v);
	assign v_w1384_v = ~(v_w1382_v & v_w1383_v);
	assign v_w14_v = ~(v_w7909_v & v_w7910_v);
	assign v_w2688_v = ~(v_w2685_v | v_w2687_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s411_v<=0;
	end
	else
	begin
	v_s411_v<=v_w462_v;
	end
	end
	assign v_w2069_v = v_w2066_v | v_w1373_v;
	assign v_w7149_v = ~(v_w7147_v | v_w7148_v);
	assign v_w7381_v = ~(v_w1846_v | v_w680_v);
	assign v_w1201_v = ~(v_w1199_v & v_w1200_v);
	assign v_w6108_v = ~(v_w6101_v & v_w6107_v);
	assign v_w6367_v = ~(v_w6365_v | v_w6366_v);
	assign v_w7126_v = ~(v_w7124_v | v_w7125_v);
	assign v_w4055_v = ~(v_w4054_v & v_s259_v);
	assign v_w7704_v = ~(v_w654_v & v_w7703_v);
	assign v_w346_v = ~(v_w7197_v & v_w7198_v);
	assign v_w3283_v = ~(v_w3279_v & v_w3282_v);
	assign v_w3211_v = ~(v_w2635_v | v_w2614_v);
	assign v_w7885_v = ~(v_s89_v & v_w7876_v);
	assign v_w6877_v = ~(v_w1788_v & v_w1126_v);
	assign v_w3204_v = ~(v_w3203_v & v_w3126_v);
	assign v_w755_v = ~(v_w813_v & v_w814_v);
	assign v_w5248_v = ~(v_w2306_v | v_w1_v);
	assign v_w7539_v = ~(v_w1188_v & v_w680_v);
	assign v_w2730_v = ~(v_w2478_v & v_w760_v);
	assign v_w449_v = ~(v_w6786_v & v_w6798_v);
	assign v_w3086_v = v_s18_v & v_w564_v;
	assign v_w3653_v = ~(v_w2459_v & v_w3652_v);
	assign v_w5081_v = v_w2460_v ^ v_w2432_v;
	assign v_w2516_v = ~(v_w558_v & v_w2327_v);
	assign v_w1772_v = ~(v_w1378_v);
	assign v_w5200_v = ~(v_w1405_v | v_w5145_v);
	assign v_w6253_v = ~(v_w657_v & v_s308_v);
	assign v_w4560_v = ~(v_w4534_v & v_w4559_v);
	assign v_w3847_v = ~(v_w2391_v & v_w3731_v);
	assign v_w1106_v = ~(v_in12_v & v_w1213_v);
	assign v_w7218_v = ~(v_s232_v & v_w7113_v);
	assign v_w5113_v = ~(v_w674_v | v_w5112_v);
	assign v_w5057_v = ~(v_w4527_v & v_w5056_v);
	assign v_w7261_v = ~(v_w7259_v | v_w7260_v);
	assign v_w2572_v = ~(v_w568_v | v_w2571_v);
	assign v_w3694_v = ~(v_w3524_v);
	assign v_w6158_v = ~(v_s236_v & v_w1528_v);
	assign v_w1130_v = ~(v_w698_v & v_s252_v);
	assign v_w2566_v = ~(v_w2560_v & v_w2565_v);
	assign v_w3224_v = ~(v_w3220_v & v_w3223_v);
	assign v_w6522_v = ~(v_w6520_v & v_w6521_v);
	assign v_w7114_v = v_s16_v & v_w7113_v;
	assign v_w151_v = v_s142_v & v_w5134_v;
	assign v_w7226_v = ~(v_s242_v & v_w7113_v);
	assign v_w5473_v = ~(v_w4863_v | v_w4712_v);
	assign v_w5776_v = ~(v_w5775_v & v_w2040_v);
	assign v_w396_v = ~(v_s509_v);
	assign v_w253_v = ~(v_w5314_v & v_w5321_v);
	assign v_w2915_v = ~(v_w2914_v | v_w993_v);
	assign v_w1231_v = ~(v_w612_v & v_s112_v);
	assign v_w6257_v = ~(v_w6029_v | v_w6256_v);
	assign v_w1324_v = ~(v_w1323_v);
	assign v_w6277_v = ~(v_w6275_v & v_w6276_v);
	assign v_w7874_v = ~(v_s197_v & v_w1993_v);
	assign v_w530_v = ~(v_w5138_v & v_w5139_v);
	assign v_w4358_v = ~(v_w8151_v);
	assign v_w1639_v = ~(v_w870_v & v_w1638_v);
	assign v_w1847_v = ~(v_w1846_v & v_w834_v);
	assign v_w2056_v = ~(v_w2009_v | v_w2055_v);
	assign v_w7468_v = ~(v_w7455_v & v_w7467_v);
	assign v_w6005_v = ~(v_w971_v ^ v_w6004_v);
	assign v_w1839_v = ~(v_w1836_v | v_w1838_v);
	assign v_w1412_v = v_w377_v ^ v_w1159_v;
	assign v_w6731_v = ~(v_w1787_v & v_w1725_v);
	assign v_w3624_v = ~(v_w3618_v & v_w3471_v);
	assign v_w2074_v = v_w2002_v & v_w1363_v;
	assign v_w4949_v = ~(v_w4941_v | v_w4589_v);
	assign v_w4528_v = ~(v_w4527_v);
	assign v_w2261_v = ~(v_w2248_v & v_w2260_v);
	assign v_w1481_v = ~(v_w666_v & v_s214_v);
	assign v_w1988_v = ~(v_w1986_v | v_w1987_v);
	assign v_w7133_v = v_w7112_v & v_s34_v;
	assign v_w6033_v = ~(v_s477_v & v_w6032_v);
	assign v_w4582_v = ~(v_w3598_v & v_w4581_v);
	assign v_w5640_v = ~(v_s203_v & v_w695_v);
	assign v_w7730_v = ~(v_s204_v & v_w7667_v);
	assign v_w7100_v = ~(v_w7098_v & v_w7099_v);
	assign v_w6106_v = ~(v_s244_v ^ v_w6105_v);
	assign v_w1261_v = ~(v_w612_v & v_s298_v);
	assign v_w7251_v = ~(v_w687_v | v_w1796_v);
	assign v_w594_v = ~(v_w1559_v & v_w1560_v);
	assign v_w1724_v = ~(v_w1052_v & v_s92_v);
	assign v_w2561_v = ~(v_w2368_v | v_w538_v);
	assign v_w6366_v = ~(v_w6018_v | v_w1465_v);
	assign v_w4453_v = ~(v_w3562_v | v_w3558_v);
	assign v_w4962_v = v_w2831_v ^ v_w4401_v;
	assign v_w2628_v = ~(v_s1_v & v_w2627_v);
	assign v_w843_v = ~(v_w705_v & v_w959_v);
	assign v_w1646_v = v_w973_v ^ v_w972_v;
	assign v_w3980_v = v_w3974_v & v_w3977_v;
	assign v_w2665_v = ~(v_w2357_v & v_s434_v);
	assign v_w6395_v = ~(v_w6383_v | v_w6394_v);
	assign v_w5906_v = ~(v_w608_v | v_w5905_v);
	assign v_w3229_v = ~(v_w3142_v | v_w2620_v);
	assign v_w8081_v = ~(v_w1923_v & v_w654_v);
	assign v_w3208_v = ~(v_w3206_v & v_w3207_v);
	assign v_w4307_v = ~(v_w4305_v | v_w4306_v);
	assign v_w3326_v = ~(v_w2815_v & v_w2634_v);
	assign v_w6843_v = ~(v_w6638_v | v_w6842_v);
	assign v_w7583_v = ~(v_w6678_v & v_w7582_v);
	assign v_w2177_v = ~(v_w701_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s157_v<=0;
	end
	else
	begin
	v_s157_v<=v_w166_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s325_v<=0;
	end
	else
	begin
	v_s325_v<=v_w351_v;
	end
	end
	assign v_w6705_v = ~(v_w656_v | v_w6704_v);
	assign v_w4562_v = ~(v_w4453_v & v_w4561_v);
	assign v_w1033_v = ~(v_w2293_v | v_w1582_v);
	assign v_w4956_v = ~(v_w4955_v & v_w673_v);
	assign v_w6828_v = ~(v_w6827_v & v_w655_v);
	assign v_w2897_v = ~(v_w2896_v);
	assign v_w1515_v = v_w1514_v | v_w1374_v;
	assign v_w3667_v = ~(v_w958_v & v_w3666_v);
	assign v_w7607_v = ~(v_w7606_v | v_w1417_v);
	assign v_w484_v = ~(v_s517_v);
	assign v_w4868_v = ~(v_w4867_v | v_w4526_v);
	assign v_w7596_v = ~(v_w961_v & v_w1902_v);
	assign v_w3122_v = ~(v_w3121_v | v_w3087_v);
	assign v_w2610_v = ~(v_w699_v & v_s211_v);
	assign v_w5607_v = ~(v_w5555_v & v_w5506_v);
	assign v_w8017_v = ~(v_w8015_v | v_w8016_v);
	assign v_w324_v = ~(v_s498_v);
	assign v_w4992_v = ~(v_w2261_v | v_w2614_v);
	assign v_w1594_v = ~(v_w1523_v | v_w1593_v);
	assign v_w7909_v = ~(v_s13_v & v_w7876_v);
	assign v_w400_v = ~(v_w3135_v & v_w3136_v);
	assign v_w5444_v = ~(v_s181_v & v_w5386_v);
	assign v_w7157_v = ~(v_w7155_v | v_w7156_v);
	assign v_w376_v = ~(v_w5832_v & v_w5839_v);
	assign v_w1913_v = ~(v_w686_v & v_w1774_v);
	assign v_w8121_v = v_w8120_v ^ v_keyinput_41_v;
	assign v_w5573_v = ~(v_w675_v & v_w5360_v);
	assign v_w526_v = ~(v_w6544_v & v_w6563_v);
	assign v_w6859_v = v_w6858_v ^ v_w1870_v;
	assign v_w4395_v = ~(v_w4393_v & v_w4394_v);
	assign v_w1468_v = ~(v_w1467_v | v_w808_v);
	assign v_w7113_v = v_w7112_v;
	assign v_w1037_v = ~(v_w1035_v & v_w1036_v);
	assign v_w7733_v = ~(v_w7660_v & v_w6917_v);
	assign v_w7761_v = ~(v_s113_v & v_w7742_v);
	assign v_w8122_v = v_w1772_v | v_w1775_v;
	assign v_w4614_v = ~(v_w674_v | v_w4613_v);
	assign v_w2879_v = ~(v_s327_v | v_w2878_v);
	assign v_w3731_v = v_w881_v;
	assign v_w2431_v = ~(v_w2428_v | v_w2430_v);
	assign v_w394_v = ~(v_w7666_v & v_w7668_v);
	assign v_w3115_v = v_w697_v & v_w3114_v;
	assign v_w5285_v = ~(v_w5283_v & v_w5284_v);
	assign v_w4693_v = ~(v_w2342_v | v_w4692_v);
	assign v_w772_v = ~(v_w1110_v | v_w1061_v);
	assign v_w3426_v = ~(v_w3424_v & v_w3425_v);
	assign v_w1730_v = ~(v_w1729_v & v_w1362_v);
	assign v_w81_v = v_s73_v & v_w7107_v;
	assign v_w4500_v = ~(v_w4452_v | v_w4499_v);
	assign v_w5470_v = ~(v_w5467_v & v_w5469_v);
	assign v_w8177_v = ~(v_w1073_v & v_w2067_v);
	assign v_w828_v = ~(v_w829_v & v_w287_v);
	assign v_w6200_v = ~(v_w6198_v | v_w6199_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s255_v<=0;
	end
	else
	begin
	v_s255_v<=v_w270_v;
	end
	end
	assign v_w4733_v = v_w820_v ^ v_w4413_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s36_v<=0;
	end
	else
	begin
	v_s36_v<=v_w43_v;
	end
	end
	assign v_w4486_v = ~(v_w958_v | v_w4485_v);
	assign v_w1510_v = ~(v_w875_v & v_s304_v);
	assign v_w2969_v = ~(v_w2966_v & v_w2968_v);
	assign v_w1375_v = ~(v_w1174_v | v_w8_v);
	assign v_w7768_v = ~(v_w6803_v | v_w1919_v);
	assign v_w2750_v = ~(v_w2749_v & v_w697_v);
	assign v_w6369_v = ~(v_w6357_v | v_w6368_v);
	assign v_w2796_v = ~(v_s476_v & v_w2776_v);
	assign v_w2808_v = ~(v_w2807_v ^ v_w581_v);
	assign v_w4111_v = ~(v_w4109_v & v_w4110_v);
	assign v_w3681_v = ~(v_w3677_v | v_w3680_v);
	assign v_w3259_v = ~(v_w810_v ^ v_w811_v);
	assign v_w7799_v = ~(v_w1734_v | v_w1782_v);
	assign v_w2160_v = ~(v_s165_v | v_w2159_v);
	assign v_w7498_v = ~(v_w7302_v & v_w7497_v);
	assign v_w5995_v = ~(v_w2117_v & v_w961_v);
	assign v_w199_v = ~(v_w5498_v & v_w5507_v);
	assign v_w8172_v = v_w6204_v | v_w6205_v;
	assign v_w1004_v = ~(v_w1289_v & v_w809_v);
	assign v_w3265_v = ~(v_w2607_v & v_w2993_v);
	assign v_w1295_v = ~(v_w1291_v | v_w1294_v);
	assign v_w6909_v = v_w1854_v & v_w1857_v;
	assign v_w8223_v = v_w2034_v & v_w903_v;
	assign v_w7119_v = ~(v_w3477_v & v_w7118_v);
	assign v_w4981_v = ~(v_w2456_v & v_w4980_v);
	assign v_w803_v = ~(v_in7_v | v_w1198_v);
	assign v_w3539_v = ~(v_w3534_v & v_w3538_v);
	assign v_w164_v = v_s155_v & v_w5134_v;
	assign v_w6989_v = ~(v_w8164_v);
	assign v_w6573_v = ~(v_w6570_v & v_w6572_v);
	assign v_w6663_v = ~(v_w6661_v & v_w758_v);
	assign v_w6468_v = ~(v_w6029_v | v_w6467_v);
	assign v_w4506_v = ~(v_w2722_v | v_w820_v);
	assign v_w3629_v = ~(v_w3628_v & v_w3593_v);
	assign v_w68_v = v_s60_v & v_w7107_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s354_v<=0;
	end
	else
	begin
	v_s354_v<=v_w392_v;
	end
	end
	assign v_w6551_v = v_w6548_v ^ v_w6550_v;
	assign v_w2461_v = ~(v_w2418_v | v_w2430_v);
	assign v_w2486_v = ~(v_w2483_v & v_w2485_v);
	assign v_w3132_v = ~(v_w8089_v);
	assign v_w7436_v = ~(v_w7375_v | v_w7378_v);
	assign v_w732_v = ~(v_s87_v & v_w1192_v);
	assign v_w1487_v = ~(v_w919_v & v_w1134_v);
	assign v_w1007_v = ~(v_w3587_v | v_w755_v);
	assign v_w1064_v = ~(v_w1300_v & v_w1301_v);
	assign v_w5235_v = ~(v_s216_v & v_w5140_v);
	assign v_w3166_v = ~(v_w3162_v | v_w3165_v);
	assign v_w6985_v = ~(v_w6978_v & v_w758_v);
	assign v_w1974_v = v_w1925_v & v_w1931_v;
	assign v_w8202_v = ~(v_w1384_v ^ v_w1999_v);
	assign v_w1700_v = v_s398_v ^ v_w1375_v;
	assign v_w511_v = ~(v_w6138_v & v_w6149_v);
	assign v_w4844_v = ~(v_w4843_v & v_w878_v);
	assign v_w853_v = ~(v_in4_v | v_w1766_v);
	assign v_w8233_v = v_w1653_v & v_w6913_v;
	assign v_w2397_v = ~(v_w2395_v | v_w2396_v);
	assign v_w6995_v = v_w1594_v ^ v_w790_v;
	assign v_w1658_v = ~(v_w1657_v);
	assign v_w7065_v = ~(v_w7063_v & v_w7064_v);
	assign v_w6814_v = ~(v_w6812_v & v_w6813_v);
	assign v_w5146_v = ~(v_w5145_v);
	assign v_w7591_v = ~(v_w7241_v | v_w7590_v);
	assign v_w1206_v = ~(v_w612_v & v_s43_v);
	assign v_w966_v = ~(v_w938_v ^ v_w965_v);
	assign v_w3958_v = ~(v_w3735_v | v_w2722_v);
	assign v_w3177_v = ~(v_w1078_v);
	assign v_w3943_v = ~(v_w3941_v | v_w3942_v);
	assign v_w7465_v = ~(v_w7449_v & v_w7452_v);
	assign v_w1392_v = ~(v_w1391_v);
	assign v_w6347_v = ~(v_s195_v & v_w888_v);
	assign v_w4773_v = v_w3177_v ^ v_w4411_v;
	assign v_w6117_v = ~(v_w1539_v ^ v_w6116_v);
	assign v_w582_v = ~(v_w585_v & v_w586_v);
	assign v_w7026_v = ~(v_w6638_v | v_w7016_v);
	assign v_w3638_v = ~(v_w3549_v & v_w3545_v);
	assign v_w7487_v = ~(v_w7485_v & v_w7486_v);
	assign v_w980_v = ~(v_w979_v);
	assign v_w7593_v = ~(v_w1996_v | v_w7592_v);
	assign v_w5522_v = ~(v_w5519_v & v_w5521_v);
	assign v_w4256_v = ~(v_w4248_v | v_w4255_v);
	assign v_w6815_v = ~(v_w6811_v | v_w6814_v);
	assign v_w4680_v = v_w3632_v ^ v_w4572_v;
	assign v_w1722_v = ~(v_w1720_v & v_w1721_v);
	assign v_w6818_v = v_s406_v & v_w656_v;
	assign v_w311_v = ~(v_w5242_v & v_w5243_v);
	assign v_w4091_v = ~(v_w4060_v & v_w4061_v);
	assign v_w4308_v = ~(v_w4299_v | v_w4307_v);
	assign v_w4418_v = ~(v_w756_v & v_w4417_v);
	assign v_w8003_v = ~(v_s280_v & v_s457_v);
	assign v_w90_v = ~(v_w7957_v & v_w7958_v);
	assign v_w8215_v = ~(v_w2745_v | v_w3050_v);
	assign v_w2599_v = ~(v_w2255_v & v_w2230_v);
	assign v_w204_v = ~(v_w5542_v & v_w5547_v);
	assign v_w2792_v = ~(v_w2484_v & v_w2791_v);
	assign v_w2544_v = ~(v_w2542_v & v_w2543_v);
	assign v_w1179_v = v_w684_v & v_s7_v;
	assign v_w930_v = ~(v_w928_v | v_w929_v);
	assign v_w115_v = ~(v_w5654_v & v_w5655_v);
	assign v_w1152_v = v_w1151_v | v_s307_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s406_v<=0;
	end
	else
	begin
	v_s406_v<=v_w455_v;
	end
	end
	assign v_w1480_v = ~(v_w1052_v & v_s215_v);
	assign v_w7156_v = v_w7113_v & v_s95_v;
	assign v_w5229_v = ~(v_w1607_v | v_w5145_v);
	assign v_w6300_v = ~(v_w6295_v ^ v_w6299_v);
	assign v_w6340_v = ~(v_w6328_v | v_w6339_v);
	assign v_w6561_v = ~(v_w6559_v | v_w6560_v);
	assign v_w5490_v = ~(v_w754_v | v_w2602_v);
	assign v_w3976_v = ~(v_w1124_v & v_w881_v);
	assign v_w2135_v = ~(v_w2124_v | v_w2134_v);
	assign v_w5693_v = ~(v_w2113_v);
	assign v_w5670_v = ~(v_s431_v & v_w695_v);
	assign v_w477_v = ~(v_w4438_v & v_w4432_v);
	assign v_w731_v = ~(v_w667_v | v_w730_v);
	assign v_w2288_v = ~(v_s476_v & v_w2287_v);
	assign v_w7597_v = ~(v_w1338_v & v_w1735_v);
	assign v_w7427_v = ~(v_w7410_v & v_w7426_v);
	assign v_w1233_v = ~(v_s161_v & v_w1192_v);
	assign v_w2847_v = ~(v_w2843_v | v_w2846_v);
	assign v_w7482_v = ~(v_w679_v | v_w1020_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s113_v<=0;
	end
	else
	begin
	v_s113_v<=v_w122_v;
	end
	end
	assign v_w4220_v = ~(v_w4206_v | v_w4219_v);
	assign v_w6504_v = ~(v_w6018_v | v_w1391_v);
	assign v_w1898_v = ~(v_w1896_v | v_w1897_v);
	assign v_w7667_v = ~(v_w654_v);
	assign v_w3520_v = v_w8246_v ^ v_keyinput_123_v;
	assign v_w1532_v = v_s285_v ^ v_s272_v;
	assign v_w6833_v = ~(v_w6831_v | v_w6832_v);
	assign v_w7515_v = ~(v_w7512_v | v_w7514_v);
	assign v_w7923_v = ~(v_s237_v & v_w6015_v);
	assign v_w6199_v = v_w1503_v & v_w6197_v;
	assign v_w4548_v = ~(v_w3639_v & v_w4547_v);
	assign v_w649_v = ~(v_w1985_v | v_w1989_v);
	assign v_w7703_v = ~(v_w7005_v & v_w7702_v);
	assign v_w1882_v = ~(v_w1815_v & v_w1881_v);
	assign v_w123_v = ~(v_w7883_v & v_w7884_v);
	assign v_w4690_v = ~(v_w4688_v | v_w4689_v);
	assign v_w2083_v = ~(v_w2080_v ^ v_w2081_v);
	assign v_w1385_v = ~(v_w1373_v | v_w1384_v);
	assign v_w4668_v = ~(v_w8248_v);
	assign v_w3069_v = ~(v_w2478_v & v_w1124_v);
	assign v_w2317_v = ~(v_w2315_v & v_w2316_v);
	assign v_w6992_v = ~(v_w6990_v & v_w6991_v);
	assign v_w3604_v = ~(v_w872_v & v_w871_v);
	assign v_w1330_v = v_s411_v ^ v_w1166_v;
	assign v_w3552_v = ~(v_w2761_v & v_w1011_v);
	assign v_w697_v = ~(v_w696_v);
	assign v_w5595_v = ~(v_w675_v & v_w5450_v);
	assign v_w2804_v = ~(v_w2478_v & v_w2803_v);
	assign v_w1277_v = ~(v_w772_v ^ v_w773_v);
	assign v_w6646_v = ~(v_w6636_v | v_w6645_v);
	assign v_w7391_v = ~(v_w687_v | v_w830_v);
	assign v_w2943_v = ~(v_w2934_v | v_w2939_v);
	assign v_w5270_v = ~(v_w5268_v | v_w5269_v);
	assign v_w2268_v = v_s249_v | v_s164_v;
	assign v_w3350_v = ~(v_w2635_v | v_w2734_v);
	assign v_w2489_v = v_s172_v & v_w604_v;
	assign v_w7059_v = ~(v_w656_v | v_w7058_v);
	assign v_w5706_v = ~(v_w5704_v | v_w5705_v);
	assign v_w2902_v = ~(v_w2478_v & v_w2901_v);
	assign v_w7385_v = ~(v_w7383_v | v_w7384_v);
	assign v_w2920_v = ~(v_w699_v & v_s351_v);
	assign v_w2043_v = ~(v_w2042_v);
	assign v_w287_v = ~(v_s494_v);
	assign v_w1359_v = ~(v_w1357_v & v_w1358_v);
	assign v_w6460_v = ~(v_w6459_v & v_w6020_v);
	assign v_w6195_v = ~(v_s226_v & v_w889_v);
	assign v_w740_v = ~(v_w1025_v & v_w784_v);
	assign v_w664_v = ~(v_w663_v | v_w2_v);
	assign v_w6060_v = ~(v_s359_v & v_w889_v);
	assign v_w7516_v = ~(v_w7279_v & v_w7515_v);
	assign v_w5671_v = ~(v_w4082_v & v_w2690_v);
	assign v_w938_v = ~(v_w8085_v);
	assign v_w5175_v = ~(v_w5146_v & v_w1329_v);
	assign v_w4533_v = ~(v_w3631_v);
	assign v_w910_v = v_w1172_v | v_w2135_v;
	assign v_w4812_v = ~(v_w4810_v | v_w4811_v);
	assign v_w2275_v = ~(v_w2273_v | v_w2274_v);
	assign v_w6962_v = ~(v_w921_v | v_w1826_v);
	assign v_w7101_v = ~(v_w1915_v | v_w6639_v);
	assign v_w4646_v = ~(v_w4645_v & v_w2341_v);
	assign v_w6875_v = ~(v_w6874_v & v_w6626_v);
	assign v_w867_v = v_w892_v & v_w893_v;
	assign v_w7866_v = ~(v_s224_v & v_w1993_v);
	assign v_w6439_v = ~(v_w6437_v & v_w6438_v);
	assign v_w1036_v = ~(v_w2272_v & v_w991_v);
	assign v_w3660_v = ~(v_w3646_v | v_w3659_v);
	assign v_w3554_v = v_w3552_v & v_w3553_v;
	assign v_w8152_v = v_w5140_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s87_v<=0;
	end
	else
	begin
	v_s87_v<=v_w95_v;
	end
	end
	assign v_w1378_v = ~(v_s100_v ^ v_w1377_v);
	assign v_w7238_v = ~(v_w7237_v | v_w6578_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s474_v<=0;
	end
	else
	begin
	v_s474_v<=v_w527_v;
	end
	end
	assign v_w4296_v = ~(v_w4295_v & v_w690_v);
	assign v_w2693_v = v_w553_v ^ v_w2692_v;
	assign v_w7838_v = ~(v_w7836_v | v_w7837_v);
	assign v_w100_v = ~(v_w7893_v & v_w7894_v);
	assign v_w7654_v = ~(v_w1979_v & v_w1972_v);
	assign v_w3105_v = ~(v_w3097_v & v_w3103_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s175_v<=0;
	end
	else
	begin
	v_s175_v<=v_w188_v;
	end
	end
	assign v_w4626_v = ~(v_w4625_v & v_w2456_v);
	assign v_w4297_v = ~(v_w2960_v | v_w4041_v);
	assign v_w7356_v = v_w7352_v | v_w7355_v;
	assign v_w1795_v = ~(v_w1758_v & v_w1794_v);
	assign v_w1831_v = ~(v_w1830_v & v_w566_v);
	assign v_w4784_v = ~(v_w4776_v & v_w4783_v);
	assign v_w8106_v = v_w939_v | v_w940_v;
	assign v_w7151_v = ~(v_w882_v | v_w529_v);
	assign v_w3936_v = ~(v_w3930_v & v_w3935_v);
	assign v_w5131_v = ~(v_w5129_v | v_w5130_v);
	assign v_w5801_v = ~(v_w892_v & v_w1119_v);
	assign v_w7263_v = ~(v_w1286_v | v_w680_v);
	assign v_w3275_v = ~(v_s292_v & v_w1_v);
	assign v_w2649_v = ~(v_w2648_v | v_w404_v);
	assign v_w7682_v = ~(v_w566_v | v_w1782_v);
	assign v_w4753_v = v_w761_v ^ v_w4412_v;
	assign v_w7627_v = ~(v_w7625_v | v_w7626_v);
	assign v_w5893_v = ~(v_w5891_v & v_w5892_v);
	assign v_w4954_v = ~(v_w4952_v | v_w4953_v);
	assign v_w2711_v = ~(v_w2484_v & v_w2706_v);
	assign v_w284_v = ~(v_w5624_v & v_w5625_v);
	assign v_w3066_v = ~(v_w3064_v & v_w3065_v);
	assign v_w919_v = ~(v_w1478_v & v_w1479_v);
	assign v_w2839_v = ~(v_w2837_v | v_w2838_v);
	assign v_w4003_v = ~(v_w4001_v & v_w4002_v);
	assign v_w8019_v = ~(v_s459_v ^ v_s295_v);
	assign v_w5666_v = ~(v_s43_v & v_w695_v);
	assign v_w279_v = ~(v_w4066_v & v_w4069_v);
	assign v_w8058_v = ~(v_w7989_v | v_w7990_v);
	assign v_w1665_v = ~(v_s336_v | v_w1464_v);
	assign v_w7327_v = ~(v_w1091_v | v_w680_v);
	assign v_w7343_v = ~(v_w687_v | v_w1678_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s205_v<=0;
	end
	else
	begin
	v_s205_v<=v_w218_v;
	end
	end
	assign v_w6278_v = v_w1610_v ^ v_w6277_v;
	assign v_w4950_v = ~(v_w4948_v | v_w4949_v);
	assign v_w5534_v = ~(v_s190_v & v_w5293_v);
	assign v_w4769_v = ~(v_w4762_v & v_w4768_v);
	assign v_w5643_v = ~(v_w420_v & v_w2910_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s223_v<=0;
	end
	else
	begin
	v_s223_v<=v_w236_v;
	end
	end
	assign v_w4376_v = ~(v_w4371_v & v_w4374_v);
	assign v_w716_v = ~(v_w999_v & v_w40_v);
	assign v_w1362_v = ~(v_w1360_v & v_w1361_v);
	assign v_w4737_v = v_w2734_v | v_w2261_v;
	assign v_w2580_v = ~(v_w2362_v | v_w314_v);
	assign v_w3201_v = ~(v_w3095_v | v_w2606_v);
	assign v_w5432_v = ~(v_w4807_v & v_w5431_v);
	assign v_w2864_v = ~(v_w2484_v & v_w2863_v);
	assign v_w1649_v = ~(v_s333_v & v_w562_v);
	assign v_w3253_v = ~(v_w2607_v & v_w2706_v);
	assign v_w6916_v = ~(v_w1657_v | v_w1651_v);
	assign v_w3506_v = ~(v_w3502_v & v_w3505_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s103_v<=0;
	end
	else
	begin
	v_s103_v<=v_w111_v;
	end
	end
	assign v_w1633_v = ~(v_w1624_v & v_w1632_v);
	assign v_w4239_v = v_w4235_v ^ v_w4238_v;
	assign v_w3509_v = ~(v_w2367_v & v_w2562_v);
	assign v_w2632_v = ~(v_w2630_v & v_w2631_v);
	assign v_w7688_v = ~(v_w7660_v & v_w7035_v);
	assign v_w2944_v = v_w2913_v | v_w2918_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s496_v<=0;
	end
	else
	begin
	v_s496_v<=v_w303_v;
	end
	end
	assign v_w2136_v = ~(v_w660_v);
	assign v_w6259_v = ~(v_w6257_v | v_w6258_v);
	assign v_w7347_v = ~(v_w7345_v | v_w7346_v);
	assign v_w553_v = ~(v_w552_v);
	assign v_w6720_v = ~(v_w6571_v | v_w1343_v);
	assign v_w1583_v = ~(v_w1576_v & v_w536_v);
	assign v_w1133_v = ~(v_w666_v & v_s225_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s371_v<=0;
	end
	else
	begin
	v_s371_v<=v_w414_v;
	end
	end
	assign v_w2312_v = v_s275_v ^ v_w2311_v;
	assign v_w1948_v = ~(v_s50_v | v_s49_v);
	assign v_w5424_v = ~(v_w4835_v & v_w5423_v);
	assign v_w5199_v = ~(v_s110_v & v_w5141_v);
	assign v_w7061_v = ~(v_w7059_v | v_w7060_v);
	assign v_w610_v = ~(v_w2025_v | v_w2026_v);
	assign v_w1541_v = ~(v_w1537_v & v_w1540_v);
	assign v_w7743_v = ~(v_s194_v & v_w7742_v);
	assign v_w94_v = ~(v_w7091_v & v_w7096_v);
	assign v_w2164_v = ~(v_w2163_v);
	assign v_w4249_v = ~(v_w2852_v & v_s329_v);
	assign v_w5119_v = ~(v_w5117_v & v_w5118_v);
	assign v_w2423_v = ~(v_w2357_v & v_s256_v);
	assign v_w6443_v = ~(v_w6400_v & v_w6398_v);
	assign v_w1504_v = ~(v_w1503_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s390_v<=0;
	end
	else
	begin
	v_s390_v<=v_w439_v;
	end
	end
	assign v_w191_v = ~(v_w5418_v & v_w5425_v);
	assign v_w7807_v = ~(v_w7805_v & v_w7806_v);
	assign v_w5395_v = ~(v_s175_v & v_w5386_v);
	assign v_w3206_v = ~(v_w2607_v & v_w2585_v);
	assign v_w7988_v = v_s468_v & v_s365_v;
	assign v_w924_v = ~(v_s326_v | v_s347_v);
	assign v_w5418_v = ~(v_s178_v & v_w5386_v);
	assign v_w4310_v = ~(v_w4054_v & v_s370_v);
	assign v_w568_v = ~(v_w2266_v & v_w2284_v);
	assign v_w7785_v = ~(v_s97_v & v_w7742_v);
	assign v_w5331_v = ~(v_w2371_v | v_w5330_v);
	assign v_w4414_v = ~(v_w3567_v & v_w4413_v);
	assign v_w579_v = ~(v_w2569_v & v_w2594_v);
	assign v_w4212_v = ~(v_w4211_v & v_w690_v);
	assign v_w3545_v = ~(v_w2991_v & v_w2980_v);
	assign v_w848_v = ~(v_in13_v | v_w1217_v);
	assign v_w6652_v = ~(v_w6648_v & v_w6651_v);
	assign v_w229_v = ~(v_w7931_v & v_w7932_v);
	assign v_w4915_v = ~(v_w4914_v & v_w673_v);
	assign v_w262_v = ~(v_w5258_v & v_w5259_v);
	assign v_w5196_v = v_s1_v & v_w2756_v;
	assign v_w8139_v = v_w8138_v ^ v_keyinput_51_v;
	assign v_w3303_v = v_w763_v ^ v_w3302_v;
	assign v_w1835_v = ~(v_w536_v);
	assign v_w997_v = ~(v_w1716_v & v_w1717_v);
	assign v_w4117_v = v_w4116_v ^ v_s281_v;
	assign v_w1196_v = ~(v_s22_v & v_w1192_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s206_v<=0;
	end
	else
	begin
	v_s206_v<=v_w219_v;
	end
	end
	assign v_w6685_v = ~(v_w1788_v & v_w1337_v);
	assign v_w3472_v = ~(v_s15_v & v_w2355_v);
	assign v_w436_v = ~(v_w916_v & v_w3202_v);
	assign v_w7082_v = v_w1838_v ^ v_w7081_v;
	assign v_w5186_v = ~(v_w5184_v | v_w5185_v);
	assign v_o2_v = v_w7980_v ^ v_w8049_v;
	assign v_w8181_v = v_w3753_v | v_w4005_v;
	assign v_w2993_v = ~(v_w2980_v);
	assign v_w892_v = v_w2117_v;
	assign v_w6358_v = ~(v_w1644_v & v_w6331_v);
	assign v_w4502_v = ~(v_w4500_v | v_w4501_v);
	assign v_w2215_v = ~(v_w2213_v & v_w2214_v);
	assign v_w353_v = ~(v_w5222_v & v_w5223_v);
	assign v_w3498_v = ~(v_w3497_v & v_w2408_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s166_v<=0;
	end
	else
	begin
	v_s166_v<=v_w175_v;
	end
	end
	assign v_w2605_v = v_w2600_v & v_w2455_v;
	assign v_w3053_v = ~(v_w699_v & v_s184_v);
	assign v_w20_v = ~(v_w7969_v & v_w7970_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s114_v<=0;
	end
	else
	begin
	v_s114_v<=v_w123_v;
	end
	end
	assign v_w2871_v = ~(v_w697_v & v_w2870_v);
	assign v_w623_v = ~(v_w3004_v | v_w3022_v);
	assign v_w7877_v = ~(v_s195_v & v_w7876_v);
	assign v_w690_v = ~(v_w688_v | v_w689_v);
	assign v_w370_v = ~(v_w5815_v & v_w5816_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s195_v<=0;
	end
	else
	begin
	v_s195_v<=v_w208_v;
	end
	end
	assign v_w2970_v = ~(v_w584_v | v_w2969_v);
	assign v_w3387_v = ~(v_w3386_v & v_w1139_v);
	assign v_w7862_v = ~(v_s234_v & v_w1993_v);
	assign v_w1380_v = ~(v_w1049_v ^ v_w1048_v);
	assign v_w4252_v = ~(v_w4250_v ^ v_w4251_v);
	assign v_w2748_v = ~(v_w2746_v & v_w2747_v);
	assign v_w8171_v = ~(v_w2380_v | v_w3503_v);
	assign v_w1922_v = ~(v_w1783_v & v_w1769_v);
	assign v_w4294_v = v_w2960_v ^ v_s364_v;
	assign v_w5925_v = ~(v_w901_v | v_w2138_v);
	assign v_w1737_v = ~(v_w1733_v | v_w1736_v);
	assign v_w6558_v = ~(v_s473_v & v_w664_v);
	assign v_w7092_v = ~(v_w656_v & v_s86_v);
	assign v_w6061_v = ~(v_w657_v & v_s86_v);
	assign v_w2362_v = ~(v_w2345_v & v_s292_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s290_v<=0;
	end
	else
	begin
	v_s290_v<=v_w310_v;
	end
	end
	assign v_w2790_v = ~(v_w558_v & v_w968_v);
	assign v_w7886_v = ~(v_w651_v & v_w7765_v);
	assign v_w5321_v = ~(v_w683_v & v_w5320_v);
	assign v_w6633_v = ~(v_w655_v & v_w6632_v);
	assign v_w2961_v = ~(v_w2960_v);
	assign v_w7377_v = ~(v_w687_v | v_w788_v);
	assign v_w5149_v = ~(v_w592_v | v_w1_v);
	assign v_w7657_v = ~(v_w2109_v & v_w2106_v);
	assign v_w4801_v = ~(v_w4799_v | v_w4800_v);
	assign v_w5054_v = v_w2337_v ^ v_w2318_v;
	assign v_w2979_v = ~(v_w2977_v & v_w2978_v);
	assign v_w5021_v = ~(v_w5019_v | v_w5020_v);
	assign v_w1267_v = ~(v_w710_v & v_s282_v);
	assign v_w6474_v = ~(v_w6473_v & v_w659_v);
	assign v_w5750_v = ~(v_w892_v & v_w567_v);
	assign v_w1298_v = ~(v_w962_v & v_w1297_v);
	assign v_w1335_v = ~(v_w1331_v | v_w1334_v);
	assign v_w6107_v = ~(v_w6106_v & v_w659_v);
	assign v_w7175_v = ~(v_w1424_v | v_w528_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s359_v<=0;
	end
	else
	begin
	v_s359_v<=v_w398_v;
	end
	end
	assign v_w2406_v = ~(v_w1131_v);
	assign v_w3849_v = ~(v_w3735_v & v_w2439_v);
	assign v_w1558_v = ~(v_w1557_v);
	assign v_w3959_v = ~(v_w881_v | v_w820_v);
	assign v_w1128_v = ~(v_w875_v & v_s288_v);
	assign v_w5391_v = ~(v_w4863_v | v_w4903_v);
	assign v_w1484_v = ~(v_s307_v ^ v_w1151_v);
	assign v_w1167_v = v_s411_v | v_w1166_v;
	assign v_w4015_v = ~(v_w3687_v & v_w4014_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s364_v<=0;
	end
	else
	begin
	v_s364_v<=v_w407_v;
	end
	end
	assign v_w2898_v = ~(v_w568_v | v_w2897_v);
	assign v_w7720_v = ~(v_w839_v | v_w1782_v);
	assign v_w3319_v = ~(v_w3314_v | v_w3318_v);
	assign v_w6280_v = ~(v_w6279_v & v_w659_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s49_v<=0;
	end
	else
	begin
	v_s49_v<=v_w57_v;
	end
	end
	assign v_w3417_v = ~(v_w3415_v | v_w3416_v);
	assign v_w7991_v = ~(v_s466_v | v_s353_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s139_v<=0;
	end
	else
	begin
	v_s139_v<=v_w148_v;
	end
	end
	assign v_w7677_v = ~(v_w7675_v | v_w7676_v);
	assign v_w8143_v = v_w8142_v ^ v_keyinput_54_v;
	assign v_w4827_v = ~(v_w878_v & v_w4558_v);
	assign v_w1163_v = v_s401_v | v_w1162_v;
	assign v_w1968_v = ~(v_w1926_v & v_w1967_v);
	assign v_w4696_v = ~(v_w2265_v & v_w851_v);
	assign v_w5182_v = ~(v_w5180_v | v_w5181_v);
	assign v_w3343_v = ~(v_w3342_v | v_w2620_v);
	assign v_w736_v = ~(v_w734_v | v_w735_v);
	assign v_w2652_v = v_w2651_v & v_s380_v;
	assign v_w2534_v = ~(v_w2525_v | v_w2533_v);
	assign v_w5895_v = ~(v_w2036_v | v_w2042_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s282_v<=0;
	end
	else
	begin
	v_s282_v<=v_w301_v;
	end
	end
	assign v_w7514_v = ~(v_w7508_v | v_w7513_v);
	assign v_w2393_v = ~(v_w699_v & v_s240_v);
	assign v_w8113_v = v_w8112_v ^ v_keyinput_36_v;
	assign v_w2779_v = ~(v_s162_v | v_w2778_v);
	assign v_w1901_v = ~(v_w1808_v | v_w1900_v);
	assign v_w6852_v = v_w656_v & v_s341_v;
	assign v_w1280_v = ~(v_w497_v ^ v_w1170_v);
	assign v_w5206_v = ~(v_w5204_v | v_w5205_v);
	assign v_w3532_v = ~(v_w2856_v | v_w2863_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s99_v<=0;
	end
	else
	begin
	v_s99_v<=v_w107_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s53_v<=0;
	end
	else
	begin
	v_s53_v<=v_w61_v;
	end
	end
	assign v_w4941_v = v_w3647_v ^ v_w4473_v;
	assign v_w3685_v = ~(v_w554_v | v_w3684_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s414_v<=0;
	end
	else
	begin
	v_s414_v<=v_w465_v;
	end
	end
	assign v_w7987_v = ~(v_s468_v | v_s365_v);
	assign v_w2818_v = ~(v_w2816_v & v_w2817_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s378_v<=0;
	end
	else
	begin
	v_s378_v<=v_w422_v;
	end
	end
	assign v_w7741_v = ~(v_w654_v & v_w7740_v);
	assign v_w638_v = v_w636_v & v_w637_v;
	assign v_w2968_v = ~(v_w2484_v & v_w2967_v);
	assign v_w5474_v = ~(v_w852_v | v_w2602_v);
	assign v_w1342_v = ~(v_w1340_v & v_w1341_v);
	assign v_w6245_v = ~(v_w6241_v ^ v_w6244_v);
	assign v_w3570_v = ~(v_w3568_v & v_w3569_v);
	assign v_w6844_v = ~(v_w6841_v | v_w6843_v);
	assign v_w2185_v = ~(v_w2169_v | v_w2184_v);
	assign v_w6129_v = ~(v_w6127_v ^ v_w6128_v);
	assign v_w7406_v = ~(v_w7404_v | v_w7405_v);
	assign v_w5134_v = ~(v_w2248_v & v_w2199_v);
	assign v_w4211_v = v_w4207_v ^ v_w4210_v;
	assign v_w7637_v = ~(v_w1796_v | v_w6585_v);
	assign v_w7222_v = ~(v_w1524_v & v_w7118_v);
	assign v_w1025_v = ~(v_in28_v & v_w1265_v);
	assign v_w6999_v = ~(v_w6998_v & v_w1915_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s203_v<=0;
	end
	else
	begin
	v_s203_v<=v_w216_v;
	end
	end
	assign v_w5280_v = ~(v_w3601_v | v_w4583_v);
	assign v_w7752_v = ~(v_w1783_v & v_w1681_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s242_v<=0;
	end
	else
	begin
	v_s242_v<=v_w255_v;
	end
	end
	assign v_w3299_v = ~(v_w3297_v | v_w3298_v);
	assign v_w717_v = ~(v_w716_v | v_s30_v);
	assign v_w8211_v = v_w8210_v ^ v_keyinput_102_v;
	assign v_w3775_v = ~(v_w3735_v | v_w2761_v);
	assign v_w2262_v = ~(v_w674_v & v_s294_v);
	assign v_w7585_v = ~(v_w7584_v & v_w1749_v);
	assign v_w4986_v = ~(v_w4979_v | v_w4985_v);
	assign v_w4749_v = ~(v_w4747_v | v_w4748_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s154_v<=0;
	end
	else
	begin
	v_s154_v<=v_w163_v;
	end
	end
	assign v_w2611_v = ~(v_w2355_v & v_s212_v);
	assign v_w1303_v = ~(v_w1302_v | v_w1180_v);
	assign v_w4572_v = ~(v_w3582_v | v_w4571_v);
	assign v_w2559_v = ~(v_w558_v & v_w2558_v);
	assign v_w1127_v = ~(v_w1520_v | v_w1522_v);
	assign v_w3331_v = ~(v_s156_v & v_w3222_v);
	assign v_w3787_v = ~(v_w3785_v | v_w3786_v);
	assign v_w1403_v = ~(v_w1401_v & v_w847_v);
	assign v_w7389_v = ~(v_w687_v | v_w944_v);
	assign v_w77_v = v_s69_v & v_w7107_v;
	assign v_w1518_v = ~(v_w666_v & v_s233_v);
	assign v_w7840_v = ~(v_w654_v & v_w7839_v);
	assign v_w5850_v = ~(v_w1521_v | v_w2135_v);
	assign v_w7975_v = ~(v_s8_v & v_w2143_v);
	assign v_w5982_v = ~(v_w5980_v & v_w5981_v);
	assign v_w2125_v = ~(v_w2109_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s295_v<=0;
	end
	else
	begin
	v_s295_v<=v_w317_v;
	end
	end
	assign v_w3688_v = ~(v_w3686_v);
	assign v_w4829_v = ~(v_w4827_v | v_w4828_v);
	assign v_w2684_v = ~(v_w2357_v & v_s427_v);
	assign v_w5452_v = ~(v_s182_v & v_w5386_v);
	assign v_w5463_v = ~(v_w2601_v & v_w820_v);
	assign v_w5455_v = ~(v_w4863_v | v_w4753_v);
	assign v_w3154_v = ~(v_w3152_v & v_w3153_v);
	assign v_w1718_v = v_s404_v ^ v_w1163_v;
	assign v_w4799_v = ~(v_w4534_v | v_w4559_v);
	assign v_w5754_v = ~(v_w5693_v | v_w5753_v);
	assign v_w4557_v = ~(v_w3549_v & v_w4556_v);
	assign v_w1148_v = v_s285_v | v_s272_v;
	assign v_w1613_v = ~(v_w1612_v);
	assign v_w3786_v = ~(v_w881_v | v_w2991_v);
	assign v_w1470_v = ~(v_s193_v & v_w562_v);
	assign v_w8186_v = v_w8185_v ^ v_keyinput_86_v;
	assign v_w6073_v = ~(v_w6071_v & v_w6072_v);
	assign v_w4309_v = ~(v_w4056_v & v_s365_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s91_v<=0;
	end
	else
	begin
	v_s91_v<=v_w99_v;
	end
	end
	assign v_w5588_v = ~(v_s116_v & v_w676_v);
	assign v_w6374_v = ~(v_s345_v ^ v_w6373_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s142_v<=0;
	end
	else
	begin
	v_s142_v<=v_w151_v;
	end
	end
	assign v_w6972_v = ~(v_w656_v | v_w6971_v);
	assign v_w6112_v = ~(v_w6087_v | v_w6091_v);
	assign v_w3790_v = ~(v_w3788_v | v_w3789_v);
	assign v_w2995_v = ~(v_w2992_v & v_w2994_v);
	assign v_w6920_v = ~(v_w6918_v & v_w6919_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s98_v<=0;
	end
	else
	begin
	v_s98_v<=v_w106_v;
	end
	end
	assign v_w3913_v = ~(v_w3801_v & v_w3912_v);
	assign v_w7228_v = ~(v_w7117_v | v_w1561_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s466_v<=0;
	end
	else
	begin
	v_s466_v<=v_w519_v;
	end
	end
	assign v_w2938_v = ~(v_w2484_v & v_w2937_v);
	assign v_w6837_v = ~(v_w1872_v ^ v_w1873_v);
	assign v_w7760_v = ~(v_w654_v & v_w7759_v);
	assign v_w4316_v = v_s369_v ^ v_w4315_v;
	assign v_w2036_v = ~(v_w2035_v | v_w1606_v);
	assign v_w76_v = v_s68_v & v_w7107_v;
	assign v_w6433_v = ~(v_w6406_v | v_w6432_v);
	assign v_w4692_v = v_w1124_v ^ v_w4415_v;
	assign v_w7532_v = ~(v_w7524_v & v_w7527_v);
	assign v_w3021_v = ~(v_w3013_v | v_w3020_v);
	assign v_w6711_v = ~(v_w1736_v ^ v_w1889_v);
	assign v_w7084_v = ~(v_w1788_v & v_w607_v);
	assign v_w4204_v = ~(v_w690_v & v_w4203_v);
	assign v_w6529_v = v_w8129_v ^ v_keyinput_46_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s318_v<=0;
	end
	else
	begin
	v_s318_v<=v_w343_v;
	end
	end
	assign v_w4394_v = ~(v_w880_v & v_w887_v);
	assign v_w8217_v = ~(v_w4697_v | v_w4698_v);
	assign v_w8248_v = v_w8247_v ^ v_keyinput_124_v;
	assign v_w4494_v = ~(v_w4492_v | v_w4493_v);
	assign v_w6070_v = ~(v_w6068_v & v_w6069_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s212_v<=0;
	end
	else
	begin
	v_s212_v<=v_w225_v;
	end
	end
	assign v_w3774_v = ~(v_w3770_v & v_w3773_v);
	assign v_w2729_v = v_w2725_v & v_w2728_v;
	assign v_w7236_v = v_s475_v | v_w1563_v;
	assign v_w3368_v = ~(v_w3366_v & v_w3367_v);
	assign v_w6601_v = ~(v_w884_v & v_w6600_v);
	assign v_w3784_v = v_w3780_v | v_w3783_v;
	assign v_w7256_v = ~(v_w7254_v & v_w7255_v);
	assign v_w2066_v = ~(v_w8203_v);
	assign v_w4882_v = ~(v_w4880_v | v_w4881_v);
	assign v_w7339_v = ~(v_w7337_v | v_w7338_v);
	assign v_w7993_v = ~(v_s465_v | v_s332_v);
	assign v_w5986_v = ~(v_w1507_v | v_w2135_v);
	assign v_w5909_v = ~(v_s158_v & v_w5786_v);
	assign v_w6262_v = ~(v_w6260_v & v_w6261_v);
	assign v_w895_v = ~(v_w1699_v);
	assign v_w564_v = v_w563_v;
	assign v_w2802_v = ~(v_w565_v & v_s216_v);
	assign v_w247_v = ~(v_w7862_v & v_w7863_v);
	assign v_w4628_v = ~(v_w4627_v & v_w878_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s164_v<=0;
	end
	else
	begin
	v_s164_v<=v_w173_v;
	end
	end
	assign v_w4357_v = ~(v_w2756_v ^ v_s389_v);
	assign v_w4811_v = ~(v_w1011_v | v_w2264_v);
	assign v_w3543_v = ~(v_w3541_v | v_w3542_v);
	assign v_w2297_v = ~(v_w2296_v);
	assign v_w5892_v = ~(v_w2117_v & v_w1853_v);
	assign v_w5184_v = ~(v_w693_v | v_w555_v);
	assign v_w1564_v = ~(v_w1563_v | v_w613_v);
	assign v_w4481_v = ~(v_w2937_v | v_w2935_v);
	assign v_w4194_v = v_w4056_v & v_s315_v;
	assign v_w7875_v = ~(v_w651_v & v_w7734_v);
	assign v_w5052_v = ~(v_w2308_v | v_w2264_v);
	assign v_w3617_v = ~(v_w3481_v | v_w3616_v);
	assign v_w328_v = ~(v_w5692_v & v_w5697_v);
	assign v_w6290_v = v_s324_v ^ v_w1626_v;
	assign v_w2110_v = ~(v_w2109_v & v_w1784_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s486_v<=0;
	end
	else
	begin
	v_s486_v<=v_w119_v;
	end
	end
	assign v_w7519_v = ~(v_w7268_v & v_w7271_v);
	assign v_w2298_v = ~(v_w2265_v & v_w2297_v);
	assign v_w2788_v = ~(v_w2774_v | v_w2787_v);
	assign v_w7372_v = ~(v_w7368_v & v_w7371_v);
	assign v_w268_v = ~(v_w5560_v & v_w5561_v);
	assign v_w2998_v = ~(v_w2990_v | v_w2997_v);
	assign v_w2664_v = ~(v_w699_v & v_s187_v);
	assign v_w266_v = ~(v_s491_v);
	assign v_w1235_v = ~(v_w1233_v & v_w1234_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s326_v<=0;
	end
	else
	begin
	v_s326_v<=v_w352_v;
	end
	end
	assign v_w466_v = ~(v_w7808_v & v_w7809_v);
	assign v_w1932_v = ~(v_w1929_v & v_w1931_v);
	assign v_w3437_v = ~(v_w3436_v & v_w3126_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s81_v<=0;
	end
	else
	begin
	v_s81_v<=v_w89_v;
	end
	end
	assign v_w6847_v = ~(v_w6845_v | v_w6846_v);
	assign v_w5297_v = ~(v_w683_v & v_w5296_v);
	assign v_w2890_v = ~(v_w2874_v);
	assign v_w3861_v = v_w2432_v ^ v_w3735_v;
	assign v_w8010_v = ~(v_w8007_v | v_w8009_v);
	assign v_w3703_v = ~(v_w3693_v | v_w3702_v);
	assign v_w4463_v = ~(v_w3648_v | v_w4462_v);
	assign v_w5267_v = ~(v_w3192_v & v_w2347_v);
	assign v_w6227_v = ~(v_w6199_v | v_w6202_v);
	assign v_w7035_v = v_w1590_v ^ v_w648_v;
	assign v_w432_v = ~(v_s514_v);
	assign v_w7407_v = ~(v_w680_v | v_w2016_v);
	assign v_w6604_v = ~(v_w6602_v | v_w6603_v);
	assign v_w2350_v = ~(v_w2282_v | v_w266_v);
	assign v_w4447_v = ~(v_w3630_v);
	assign v_w1076_v = ~(v_w3037_v & v_w3038_v);
	assign v_w3234_v = ~(v_w820_v & v_w2639_v);
	assign v_w3782_v = ~(v_w967_v | v_w3735_v);
	assign v_w6415_v = ~(v_s122_v & v_w6387_v);
	assign v_w1632_v = ~(v_w1630_v & v_w1631_v);
	assign v_w2427_v = ~(v_w2419_v & v_w2426_v);
	assign v_w6883_v = ~(v_w6571_v | v_w1674_v);
	assign v_w4306_v = ~(v_w4300_v | v_w4303_v);
	assign v_w5181_v = v_w5141_v & v_s82_v;
	assign v_w2812_v = ~(v_w2355_v & v_s210_v);
	assign v_w7774_v = ~(v_w1075_v | v_w1782_v);
	assign v_w6263_v = v_w1610_v ^ v_w6262_v;
	assign v_w3390_v = ~(v_w2635_v | v_w2906_v);
	assign v_w3369_v = ~(v_w3077_v);
	assign v_w6610_v = ~(v_w6609_v & v_w655_v);
	assign v_w5755_v = ~(v_s272_v | v_w2135_v);
	assign v_w3161_v = ~(v_w3109_v & v_w2439_v);
	assign v_w7545_v = ~(v_w7248_v | v_w7244_v);
	assign v_w5574_v = ~(v_s210_v & v_w676_v);
	assign v_w3345_v = ~(v_w2745_v | v_w3049_v);
	assign v_w4599_v = v_w3098_v ^ v_w4419_v;
	assign v_w1920_v = ~(v_w1000_v | v_w1919_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s337_v<=0;
	end
	else
	begin
	v_s337_v<=v_w368_v;
	end
	end
	assign v_w321_v = ~(v_w5011_v & v_w5012_v);
	assign v_w558_v = ~(v_w557_v);
	assign v_w5249_v = v_w5140_v & v_s237_v;
	assign v_w3585_v = ~(v_w3576_v | v_w3584_v);
	assign v_w5701_v = ~(v_w1188_v | v_w2138_v);
	assign v_w5511_v = ~(v_w5509_v & v_w5510_v);
	assign v_w2450_v = ~(v_w2446_v & v_w2449_v);
	assign v_w6213_v = ~(v_w6212_v ^ v_s224_v);
	assign v_w7174_v = ~(v_s373_v & v_w7113_v);
	assign v_w2178_v = ~(v_w947_v);
	assign v_w2318_v = ~(v_w2317_v);
	assign v_w7045_v = ~(v_w1842_v ^ v_w1548_v);
	assign v_w3191_v = ~(v_w3186_v ^ v_w966_v);
	assign v_w8013_v = ~(v_w8005_v & v_w8012_v);
	assign v_w6493_v = ~(v_w6491_v & v_w6492_v);
	assign v_w6211_v = ~(v_w6209_v & v_w6210_v);
	assign v_w7581_v = ~(v_w7579_v & v_w7580_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s193_v<=0;
	end
	else
	begin
	v_s193_v<=v_w206_v;
	end
	end
	assign v_w5145_v = ~(v_w1192_v & v_w693_v);
	assign v_w7681_v = ~(v_w7047_v | v_w1919_v);
	assign v_w7797_v = ~(v_s80_v & v_w7742_v);
	assign v_w4068_v = v_w4067_v ^ v_w4044_v;
	assign v_w453_v = ~(v_w5914_v & v_w5921_v);
	assign v_w1478_v = ~(v_w1475_v | v_w1477_v);
	assign v_w1141_v = ~(v_w1985_v | v_w6576_v);
	assign v_w4168_v = ~(v_w4166_v | v_w4167_v);
	assign v_w7191_v = ~(v_w1644_v | v_w529_v);
	assign v_w8127_v = v_w6713_v | v_w1919_v;
	assign v_w6091_v = ~(v_w1557_v ^ v_w6090_v);
	assign v_w3749_v = v_w3745_v | v_w3748_v;
	assign v_w5049_v = ~(v_w674_v & v_s281_v);
	assign v_w2948_v = v_w2942_v & v_w2947_v;
	assign v_w96_v = ~(v_w7766_v & v_w7767_v);
	assign v_o1_v = ~(v_w8051_v ^ v_w8052_v);
	assign v_w5867_v = ~(v_w5865_v & v_w5866_v);
	assign v_w2682_v = ~(v_w2478_v & v_w755_v);
	assign v_w2922_v = v_w387_v ^ v_w2644_v;
	assign v_w1746_v = ~(v_w1326_v | v_w1745_v);
	assign v_w5806_v = ~(v_w1820_v | v_w2138_v);
	assign v_w5169_v = v_w5141_v & v_s32_v;
	assign v_w74_v = v_s66_v & v_w7107_v;
	assign v_w1523_v = ~(v_w834_v | v_w1026_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s370_v<=0;
	end
	else
	begin
	v_s370_v<=v_w413_v;
	end
	end
	assign v_w2625_v = ~(v_w2624_v | v_w1138_v);
	assign v_w1994_v = ~(v_s10_v & v_w1993_v);
	assign v_w5485_v = ~(v_w5484_v | v_w4688_v);
	assign v_w7005_v = ~(v_w7001_v | v_w7004_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s467_v<=0;
	end
	else
	begin
	v_s467_v<=v_w520_v;
	end
	end
	assign v_w992_v = ~(v_w2341_v | v_w616_v);
	assign v_w5245_v = ~(v_w5145_v | v_w1517_v);
	assign v_w580_v = ~(v_w2587_v & v_w2593_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s305_v<=0;
	end
	else
	begin
	v_s305_v<=v_w328_v;
	end
	end
	assign v_w5917_v = ~(v_w5916_v & v_w2113_v);
	assign v_w1070_v = ~(v_w1405_v | v_w808_v);
	assign v_w2496_v = ~(v_w604_v & v_s258_v);
	assign v_w2775_v = v_w711_v & v_w2147_v;
	assign v_w1771_v = ~(v_w8_v | v_w1770_v);
	assign v_w3116_v = ~(v_w3112_v | v_w3115_v);
	assign v_w3956_v = ~(v_w3951_v & v_w3955_v);
	assign v_w7740_v = ~(v_w6903_v & v_w7739_v);
	assign v_w1162_v = v_w1161_v | v_s399_v;
	assign v_w2225_v = ~(v_w2223_v & v_w2224_v);
	assign v_w3443_v = ~(v_w2991_v & v_w2639_v);
	assign v_w6187_v = v_s226_v ^ v_w1503_v;
	assign v_w47_v = ~(v_w4037_v | v_w4038_v);
	assign v_w7602_v = ~(v_w7601_v & v_w1679_v);
	assign v_w2477_v = ~(v_w2453_v & v_w2476_v);
	assign v_w7633_v = ~(v_w6586_v | v_w7632_v);
	assign v_w412_v = ~(v_w4842_v & v_w4857_v);
	assign v_w6533_v = ~(v_w5969_v & v_w6532_v);
	assign v_w3370_v = v_w8237_v ^ v_keyinput_118_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s481_v<=0;
	end
	else
	begin
	v_s481_v<=v_w27_v;
	end
	end
	assign v_w719_v = v_w909_v & v_w363_v;
	assign v_w6170_v = ~(v_w657_v & v_s288_v);
	assign v_w7023_v = ~(v_w7021_v & v_w7022_v);
	assign v_w297_v = ~(v_w3311_v & v_w3319_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s161_v<=0;
	end
	else
	begin
	v_s161_v<=v_w170_v;
	end
	end
	assign v_w7404_v = ~(v_w687_v | v_w596_v);
	assign v_w6802_v = ~(v_w928_v | v_w1818_v);
	assign v_w8090_v = v_w2926_v | v_w2620_v;
	assign v_w8112_v = ~(v_w2258_v & v_w2259_v);
	assign v_w5527_v = v_w8176_v ^ v_keyinput_80_v;
	assign v_w1567_v = ~(v_w1565_v & v_w1566_v);
	assign v_w2720_v = ~(v_w2717_v | v_w2719_v);
	assign v_w4914_v = ~(v_w4907_v & v_w4913_v);
	assign v_w2247_v = ~(v_s1_v & v_w2246_v);
	assign v_w1492_v = ~(v_w562_v & v_s222_v);
	assign v_w2017_v = ~(v_w2016_v ^ v_w1999_v);
	assign v_w7370_v = ~(v_w687_v | v_w1100_v);
	assign v_w845_v = ~(v_w1386_v | v_w808_v);
	assign v_w6124_v = ~(v_w5876_v & v_w6123_v);
	assign v_w7230_v = ~(v_s267_v & v_w7113_v);
	assign v_w1867_v = ~(v_w1678_v & v_w1866_v);
	assign v_w1938_v = ~(v_w1936_v & v_w1937_v);
	assign v_w3325_v = ~(v_w2831_v & v_w2639_v);
	assign v_w1930_v = ~(v_w8_v | v_w1178_v);
	assign v_w2022_v = v_w575_v ^ v_w2019_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s140_v<=0;
	end
	else
	begin
	v_s140_v<=v_w149_v;
	end
	end
	assign v_w4093_v = ~(v_w4089_v & v_w4092_v);
	assign v_w3026_v = ~(v_w2484_v & v_w3025_v);
	assign v_w1533_v = ~(v_w1532_v | v_w1180_v);
	assign v_w1833_v = ~(v_w575_v | v_w536_v);
	assign v_w4965_v = v_w3646_v ^ v_w4470_v;
	assign v_w5217_v = ~(v_w1467_v | v_w5145_v);
	assign v_w4973_v = ~(v_w4966_v & v_w4972_v);
	assign v_w802_v = ~(v_w800_v & v_w801_v);
	assign v_w2203_v = ~(v_w2201_v & v_w2202_v);
	assign v_w3145_v = ~(v_w3138_v & v_w3144_v);
	assign v_w1678_v = ~(v_w1676_v & v_w1677_v);
	assign v_w1785_v = ~(v_w1778_v & v_w1784_v);
	assign v_w2980_v = ~(v_w2975_v | v_w2979_v);
	assign v_w3059_v = ~(v_w593_v & v_s77_v);
	assign v_w8207_v = v_w8206_v ^ v_keyinput_99_v;
	assign v_w4658_v = ~(v_w2448_v & v_w3077_v);
	assign v_w1081_v = ~(v_w2982_v & v_w2986_v);
	assign v_w3664_v = ~(v_w3640_v | v_w3663_v);
	assign v_w7459_v = ~(v_w7457_v & v_w7458_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s214_v<=0;
	end
	else
	begin
	v_s214_v<=v_w227_v;
	end
	end
	assign v_w1894_v = ~(v_w1891_v);
	assign v_w5955_v = ~(v_w2051_v ^ v_w5954_v);
	assign v_w7280_v = ~(v_w680_v | v_w1119_v);
	assign v_w8146_v = v_w974_v ^ v_w975_v;
	assign v_w2623_v = ~(v_w8194_v);
	assign v_w7250_v = ~(v_w6586_v | v_w680_v);
	assign v_w8242_v = ~(v_w3017_v | v_w4041_v);
	assign v_w2874_v = ~(v_w2869_v | v_w2873_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s278_v<=0;
	end
	else
	begin
	v_s278_v<=v_w297_v;
	end
	end
	assign v_w4597_v = ~(v_w3087_v | v_w2264_v);
	assign v_w3019_v = ~(v_w3018_v & v_w569_v);
	assign v_w7396_v = ~(v_w680_v | v_w567_v);
	assign v_w2309_v = ~(v_w2308_v);
	assign v_w7680_v = ~(v_s245_v & v_w7667_v);
	assign v_w2420_v = ~(v_s156_v & v_w697_v);
	assign v_w7379_v = ~(v_w7375_v & v_w7378_v);
	assign v_w2030_v = ~(v_w766_v ^ v_w722_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s167_v<=0;
	end
	else
	begin
	v_s167_v<=v_w177_v;
	end
	end
	assign v_w101_v = ~(v_w7955_v & v_w7956_v);
	assign v_w889_v = ~(v_w891_v ^ v_w34_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s475_v<=0;
	end
	else
	begin
	v_s475_v<=v_w528_v;
	end
	end
	assign v_w6693_v = ~(v_w6691_v & v_w6692_v);
	assign v_w4526_v = ~(v_w4525_v);
	assign v_w5030_v = ~(v_w5028_v & v_w5029_v);
	assign v_w7529_v = ~(v_w7521_v | v_w7528_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s25_v<=0;
	end
	else
	begin
	v_s25_v<=v_w27_v;
	end
	end
	assign v_w7358_v = ~(v_w680_v | v_w1650_v);
	assign v_w6959_v = ~(v_w6954_v | v_w6958_v);
	assign v_w4793_v = ~(v_w4791_v | v_w4792_v);
	assign v_w5352_v = ~(v_w5003_v & v_w5351_v);
	assign v_w1770_v = v_w778_v & v_w1177_v;
	assign v_w1742_v = ~(v_w1741_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s28_v<=0;
	end
	else
	begin
	v_s28_v<=v_w31_v;
	end
	end
	assign v_w3195_v = ~(v_w3193_v & v_w3194_v);
	assign v_w1200_v = ~(v_w612_v & v_s431_v);
	assign v_w3531_v = ~(v_w2916_v | v_w2910_v);
	assign v_w5495_v = ~(v_w5493_v | v_w5494_v);
	assign v_w7227_v = ~(v_w1557_v | v_w528_v);
	assign v_w2875_v = ~(v_w2874_v | v_w538_v);
	assign v_w916_v = v_w914_v & v_w915_v;
	assign v_w6309_v = ~(v_w5738_v & v_w6308_v);
	assign v_w1220_v = ~(v_w1218_v & v_w1219_v);
	assign v_w1826_v = ~(v_w1135_v | v_w919_v);
	assign v_w1028_v = v_w1026_v ^ v_w1027_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s380_v<=0;
	end
	else
	begin
	v_s380_v<=v_w426_v;
	end
	end
	assign v_w4288_v = ~(v_w4286_v & v_w4287_v);
	assign v_w3851_v = ~(v_w3849_v & v_w3850_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s367_v<=0;
	end
	else
	begin
	v_s367_v<=v_w410_v;
	end
	end
	assign v_w1885_v = ~(v_w1726_v & v_w998_v);
	assign v_w1544_v = ~(v_w874_v & v_s273_v);
	assign v_w1803_v = ~(v_w893_v);
	assign v_w5777_v = ~(v_w2044_v & v_w2033_v);
	assign v_w4344_v = ~(v_w4342_v | v_w4343_v);
	assign v_w17_v = ~(v_w5680_v & v_w5681_v);
	assign v_w461_v = ~(v_s516_v);
	assign v_w5730_v = ~(v_w5724_v & v_w5729_v);
	assign v_w7441_v = ~(v_w687_v | v_w1606_v);
	assign v_w3864_v = ~(v_w881_v | v_w2317_v);
	assign v_o22_v = ~(v_s474_v ^ v_s376_v);
	assign v_w4694_v = ~(v_w4691_v | v_w4693_v);
	assign v_w2787_v = ~(v_w967_v | v_w617_v);
	assign v_w6205_v = ~(v_w6018_v | v_w1503_v);
	assign v_w6754_v = ~(v_w6750_v | v_w6753_v);
	assign v_w4379_v = ~(v_w4370_v | v_w4378_v);
	assign v_w4529_v = ~(v_w4524_v | v_w4528_v);
	assign v_w7588_v = ~(v_w934_v | v_w7587_v);
	assign v_w2370_v = ~(v_w2369_v);
	assign v_w1748_v = ~(v_w1310_v | v_w1747_v);
	assign v_w3503_v = ~(v_w2562_v | v_w2367_v);
	assign v_w7642_v = ~(v_w1913_v | v_w7641_v);
	assign v_w5213_v = ~(v_w8205_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s117_v<=0;
	end
	else
	begin
	v_s117_v<=v_w126_v;
	end
	end
	assign v_w2004_v = ~(v_w1999_v ^ v_w998_v);
	assign v_w797_v = ~(v_w997_v | v_w1726_v);
	assign v_w1091_v = ~(v_w1089_v | v_w1090_v);
	assign v_w7747_v = ~(v_w6880_v & v_w7746_v);
	assign v_w215_v = ~(v_w5576_v & v_w5577_v);
	assign v_w365_v = ~(v_s503_v);
	assign v_w4756_v = ~(v_w674_v & v_s394_v);
	assign v_w5736_v = ~(v_w1642_v | v_w2138_v);
	assign v_w4112_v = v_w4108_v ^ v_w4111_v;
	assign v_w4349_v = ~(v_w4346_v ^ v_w4348_v);
	assign v_w6739_v = ~(v_w6637_v | v_w6735_v);
	assign v_w2607_v = ~(v_w2606_v);
	assign v_w3542_v = ~(v_w2874_v | v_w1017_v);
	assign v_w783_v = v_in28_v ^ v_w1265_v;
	assign v_w6738_v = ~(v_w8080_v);
	assign v_w7063_v = ~(v_w656_v & v_s271_v);
	assign v_w3815_v = v_w3811_v | v_w3814_v;
	assign v_w7171_v = ~(v_w6457_v | v_w529_v);
	assign v_w7533_v = ~(v_w7531_v & v_w7532_v);
	assign v_w7355_v = ~(v_w7353_v | v_w7354_v);
	assign v_w3186_v = ~(v_w3185_v & v_w3104_v);
	assign v_w1561_v = ~(v_w744_v ^ v_w704_v);
	assign v_w557_v = ~(v_w537_v);
	assign v_w1527_v = v_w828_v & v_s7_v;
	assign v_w7180_v = ~(v_w1443_v | v_w7117_v);
	assign v_w7934_v = ~(v_w527_v & v_w1606_v);
	assign v_w6597_v = ~(v_w936_v);
	assign v_w8241_v = v_w8240_v ^ v_keyinput_120_v;
	assign v_w4922_v = ~(v_w4921_v & v_w878_v);
	assign v_w4101_v = v_s241_v ^ v_w2312_v;
	assign v_w6435_v = ~(v_w657_v & v_s354_v);
	assign v_w864_v = ~(v_w862_v | v_w863_v);
	assign v_w7048_v = ~(v_w7047_v);
	assign v_w6109_v = ~(v_w6018_v | v_w1539_v);
	assign v_w2058_v = ~(v_w1999_v ^ v_w1091_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s285_v<=0;
	end
	else
	begin
	v_s285_v<=v_w305_v;
	end
	end
	assign v_w3393_v = ~(v_w3109_v & v_w2399_v);
	assign v_w6361_v = v_s344_v ^ v_w1465_v;
	assign v_w5997_v = ~(v_w1290_v | v_w2135_v);
	assign v_w7196_v = ~(v_w7117_v | v_w1628_v);
	assign v_w6450_v = ~(v_w6018_v | v_w1424_v);
	assign v_w2701_v = ~(v_w2699_v & v_w2700_v);
	assign v_w3867_v = ~(v_w2318_v | v_w3735_v);
	assign v_w7336_v = ~(v_w7334_v | v_w7335_v);
	assign v_w4687_v = ~(v_w4684_v | v_w4686_v);
	assign v_w2402_v = ~(v_s261_v & v_w697_v);
	assign v_w5791_v = ~(v_w2021_v ^ v_w2022_v);
	assign v_w3138_v = ~(v_w3137_v & v_w3126_v);
	assign v_w6612_v = ~(v_w6592_v & v_w893_v);
	assign v_w7729_v = ~(v_w654_v & v_w7728_v);
	assign v_w221_v = ~(v_w7933_v & v_w7934_v);
	assign v_w5371_v = ~(v_w4941_v | v_w5123_v);
	assign v_w7904_v = ~(v_w651_v & v_w7820_v);
	assign v_w492_v = ~(v_w5992_v & v_w5998_v);
	assign v_w2835_v = ~(v_w2832_v & v_w2834_v);
	assign v_w2226_v = ~(v_w2222_v | v_w2225_v);
	assign v_w6986_v = ~(v_w6984_v & v_w6985_v);
	assign v_w4865_v = ~(v_w4863_v | v_w4864_v);
	assign v_w5660_v = ~(v_s95_v & v_w695_v);
	assign v_w787_v = ~(v_w1996_v | v_w1980_v);
	assign v_w5205_v = ~(v_w5145_v | v_w1427_v);
	assign v_w7664_v = ~(v_w7662_v | v_w7663_v);
	assign v_w7383_v = ~(v_w680_v | v_w1027_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s355_v<=0;
	end
	else
	begin
	v_s355_v<=v_w393_v;
	end
	end
	assign v_w6194_v = ~(v_w6180_v | v_w6193_v);
	assign v_w2460_v = ~(v_w2409_v);
	assign v_w6294_v = ~(v_w6268_v | v_w6272_v);
	assign v_w7408_v = ~(v_w687_v | v_w602_v);
	assign v_w631_v = v_w629_v & v_w630_v;
	assign v_w1672_v = ~(v_w875_v & v_s345_v);
	assign v_w1818_v = ~(v_w1401_v | v_w1817_v);
	assign v_w3495_v = ~(v_w2419_v | v_w2426_v);
	assign v_w7860_v = ~(v_s236_v & v_w1993_v);
	assign v_o19_v = v_s455_v ^ v_w8053_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s116_v<=0;
	end
	else
	begin
	v_s116_v<=v_w125_v;
	end
	end
	assign v_w3084_v = ~(v_w2681_v | v_w941_v);
	assign v_w2896_v = v_s327_v ^ v_w2878_v;
	assign v_w3603_v = ~(v_w3597_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s454_v<=0;
	end
	else
	begin
	v_s454_v<=v_w507_v;
	end
	end
	assign v_w7955_v = ~(v_s93_v & v_w2143_v);
	assign v_w6201_v = ~(v_w6168_v & v_w6173_v);
	assign v_w2344_v = ~(v_w2340_v & v_w2343_v);
	assign v_w2054_v = ~(v_w723_v ^ v_w1096_v);
	assign v_w4416_v = ~(v_w3574_v & v_w4415_v);
	assign v_w5642_v = ~(v_s333_v & v_w695_v);
	assign v_w781_v = ~(v_w3568_v & v_w3579_v);
	assign v_w2045_v = v_w2043_v & v_w2044_v;
	assign v_w5882_v = v_w8148_v ^ v_keyinput_58_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s294_v<=0;
	end
	else
	begin
	v_s294_v<=v_w316_v;
	end
	end
	assign v_w1234_v = ~(v_w612_v & v_s366_v);
	assign v_w3622_v = ~(v_w3621_v & v_w555_v);
	assign v_w547_v = v_s395_v | v_s473_v;
	assign v_w4948_v = ~(v_w4946_v | v_w4947_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s85_v<=0;
	end
	else
	begin
	v_s85_v<=v_w93_v;
	end
	end
	assign v_w1673_v = ~(v_w1671_v & v_w1672_v);
	assign v_w7894_v = ~(v_w651_v & v_w7789_v);
	assign v_w6269_v = ~(v_s207_v & v_w888_v);
	assign v_w1765_v = ~(v_w612_v & v_s20_v);
	assign v_w2062_v = v_w1401_v & v_w2007_v;
	assign v_w2421_v = ~(v_s258_v & v_w593_v);
	assign v_w8175_v = v_w3685_v | v_w4027_v;
	assign v_w3429_v = ~(v_w2681_v | v_w939_v);
	assign v_w6938_v = ~(v_w656_v | v_w6937_v);
	assign v_w4023_v = ~(v_w2241_v & v_w4020_v);
	assign v_w7724_v = ~(v_s206_v & v_w7667_v);
	assign v_w836_v = ~(v_w1491_v & v_w1492_v);
	assign v_w3841_v = ~(v_w2558_v & v_w3731_v);
	assign v_w5864_v = ~(v_w5862_v | v_w5863_v);
	assign v_w4189_v = ~(v_w4187_v & v_w4188_v);
	assign v_w4401_v = ~(v_w2803_v | v_w4400_v);
	assign v_w5407_v = ~(v_w4876_v | v_w5406_v);
	assign v_w4007_v = ~(v_w3750_v & v_w4006_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s18_v<=0;
	end
	else
	begin
	v_s18_v<=v_w20_v;
	end
	end
	assign v_w2800_v = ~(v_w2799_v | v_w568_v);
	assign v_w6660_v = v_w1746_v ^ v_w6659_v;
	assign v_w132_v = ~(v_w7941_v & v_w7942_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s30_v<=0;
	end
	else
	begin
	v_s30_v<=v_w33_v;
	end
	end
	assign v_w3739_v = ~(v_w3199_v | v_w3731_v);
	assign v_w195_v = ~(v_w5452_v & v_w5461_v);
	assign v_w585_v = ~(v_w2894_v & v_w638_v);
	assign v_w5904_v = ~(v_w5902_v & v_w5903_v);
	assign v_w230_v = ~(v_w5234_v & v_w5235_v);
	assign v_w5029_v = ~(v_w2265_v & v_w2558_v);
	assign v_w263_v = ~(v_s490_v);
	assign v_w5480_v = ~(v_s185_v & v_w5386_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s276_v<=0;
	end
	else
	begin
	v_s276_v<=v_w294_v;
	end
	end
	assign v_w5233_v = ~(v_w2799_v | v_w1_v);
	assign v_w4134_v = ~(v_w4088_v | v_w4133_v);
	assign v_w3300_v = ~(v_w2607_v & v_w3077_v);
	assign v_w3430_v = v_w940_v ^ v_w3429_v;
	assign v_w6702_v = ~(v_w6695_v & v_w6701_v);
	assign v_w2999_v = ~(v_w2789_v ^ v_w2793_v);
	assign v_w1900_v = ~(v_w1809_v | v_w1899_v);
	assign v_w2842_v = ~(v_s202_v & v_w2355_v);
	assign v_w288_v = ~(v_w5964_v & v_w5965_v);
	assign v_w3594_v = v_w3592_v & v_w3593_v;
	assign v_w4669_v = ~(v_w4667_v | v_w4668_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s504_v<=0;
	end
	else
	begin
	v_s504_v<=v_w366_v;
	end
	end
	assign v_w7580_v = ~(v_w1741_v | v_w1887_v);
	assign v_w8092_v = v_w8091_v ^ v_keyinput_20_v;
	assign v_w281_v = ~(v_w5622_v & v_w5623_v);
	assign v_w3271_v = ~(v_w2766_v & v_w2634_v);
	assign v_w5031_v = v_w2562_v ^ v_w4398_v;
	assign v_w745_v = ~(v_w744_v & v_w704_v);
	assign v_w7488_v = ~(v_w7484_v & v_w7487_v);
	assign v_w4409_v = ~(v_w968_v | v_w4408_v);
	assign v_w3521_v = ~(v_w2803_v);
	assign v_w5891_v = ~(v_w662_v & v_w1135_v);
	assign v_w3464_v = v_w3456_v ^ v_w3463_v;
	assign v_w460_v = ~(v_w5943_v & v_w5944_v);
	assign v_w5117_v = ~(v_w674_v & v_s256_v);
	assign v_w5059_v = v_s279_v & v_w674_v;
	assign v_w7384_v = ~(v_w687_v | v_w1026_v);
	assign v_w6736_v = ~(v_w6638_v | v_w6735_v);
	assign v_w1058_v = ~(v_in8_v ^ v_w1201_v);
	assign v_w2099_v = ~(v_w2096_v & v_w2098_v);
	assign v_w7466_v = ~(v_w7446_v | v_w7465_v);
	assign v_w4120_v = ~(v_w4118_v & v_w4119_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s270_v<=0;
	end
	else
	begin
	v_s270_v<=v_w288_v;
	end
	end
	assign v_w3541_v = ~(v_w956_v);
	assign v_w1841_v = ~(v_w603_v & v_w1840_v);
	assign v_w5434_v = ~(v_s180_v & v_w5386_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s100_v<=0;
	end
	else
	begin
	v_s100_v<=v_w108_v;
	end
	end
	assign v_w5913_v = ~(v_w1363_v | v_w2138_v);
	assign v_w3242_v = ~(v_w3238_v | v_w3241_v);
	assign v_w3866_v = ~(v_w2400_v | v_w3731_v);
	assign v_w1820_v = ~(v_w1678_v);
	assign v_w3465_v = v_w710_v | v_w3464_v;
	assign v_w1409_v = ~(v_w666_v & v_s88_v);
	assign v_w8220_v = v_w8219_v ^ v_keyinput_107_v;
	assign v_w5_v = ~(v_w5618_v & v_w5619_v);
	assign v_w470_v = ~(v_w7846_v & v_w7847_v);
	assign v_w3433_v = ~(v_w3431_v & v_w3432_v);
	assign v_w970_v = v_w2056_v | v_w2057_v;
	assign v_w5204_v = ~(v_w693_v | v_w2984_v);
	assign v_w4573_v = ~(v_w3632_v);
	assign v_w6156_v = ~(v_w6155_v ^ v_s288_v);
	assign v_w1463_v = ~(v_s334_v | v_w1462_v);
	assign v_w5766_v = ~(v_w2067_v & v_w2069_v);
	assign v_w2202_v = ~(v_s145_v | v_s144_v);
	assign v_w7868_v = ~(v_s215_v & v_w1993_v);
	assign v_w7712_v = ~(v_s223_v & v_w7667_v);
	assign v_w1854_v = ~(v_w1606_v & v_w1853_v);
	assign v_w3077_v = ~(v_w3075_v & v_w3076_v);
	assign v_w6698_v = ~(v_w6696_v & v_w6697_v);
	assign v_w737_v = ~(v_w8083_v);
	assign v_w7903_v = ~(v_s26_v & v_w1993_v);
	assign v_w2755_v = ~(v_s110_v & v_w564_v);
	assign v_w3147_v = ~(v_w3145_v | v_w3146_v);
	assign v_w2155_v = ~(v_w2154_v);
	assign v_w5798_v = ~(v_w2074_v | v_w2003_v);
	assign v_w967_v = ~(v_w1084_v | v_w1085_v);
	assign v_w2337_v = ~(v_w2327_v | v_w2336_v);
	assign v_w7502_v = ~(v_w7294_v | v_w7501_v);
	assign v_w6626_v = ~(v_w6602_v);
	assign v_w7573_v = ~(v_w7572_v & v_w6870_v);
	assign v_w7666_v = ~(v_w654_v & v_w7665_v);
	assign v_w2827_v = ~(v_w2825_v | v_w2826_v);
	assign v_w7095_v = ~(v_w536_v | v_w6579_v);
	assign v_w699_v = v_w698_v;
	assign v_w2675_v = ~(v_w558_v & v_w871_v);
	assign v_w4295_v = ~(v_w4293_v ^ v_w4294_v);
	assign v_w409_v = ~(v_w5648_v & v_w5649_v);
	assign v_w2073_v = ~(v_w2003_v | v_w2072_v);
	assign v_w4199_v = v_w4190_v ^ v_s314_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s72_v<=0;
	end
	else
	begin
	v_s72_v<=v_w80_v;
	end
	end
	assign v_w2951_v = ~(v_w2949_v & v_w2950_v);
	assign v_w7_v = ~(v_w7110_v & v_w7111_v);
	assign v_w2811_v = ~(v_w2809_v & v_w2810_v);
	assign v_w209_v = ~(v_w7735_v & v_w7736_v);
	assign v_w7322_v = ~(v_w680_v | v_w1817_v);
	assign v_w5064_v = ~(v_w2407_v & v_w5063_v);
	assign v_w4886_v = ~(v_w2342_v | v_w4885_v);
	assign v_w4826_v = ~(v_w4825_v & v_w2341_v);
	assign v_w7155_v = ~(v_w1775_v | v_w529_v);
	assign v_w4164_v = v_w4160_v ^ v_w4163_v;
	assign v_w5783_v = ~(v_w662_v & v_w607_v);
	assign v_w3334_v = ~(v_w3121_v | v_w2335_v);
	assign v_w5125_v = ~(v_w5124_v | v_w4588_v);
	assign v_w5933_v = ~(v_w5931_v | v_w5932_v);
	assign v_w3471_v = ~(v_w3470_v);
	assign v_w4511_v = ~(v_w3077_v | v_w1124_v);
	assign v_w7973_v = ~(v_s11_v & v_w2143_v);
	assign v_w4601_v = ~(v_w2448_v & v_w2671_v);
	assign v_w3652_v = ~(v_w3495_v | v_w2409_v);
	assign v_w381_v = ~(v_w7939_v & v_w7940_v);
	assign v_w6351_v = v_w1465_v & v_w6349_v;
	assign v_w2742_v = ~(v_w558_v & v_w760_v);
	assign v_w2359_v = ~(v_w2358_v & v_s296_v);
	assign v_w382_v = ~(v_w5218_v & v_w5219_v);
	assign v_w4591_v = ~(v_w4587_v | v_w4590_v);
	assign v_w6518_v = ~(v_w6019_v | v_w6517_v);
	assign v_w886_v = ~(v_w2284_v & v_w4040_v);
	assign v_w2149_v = ~(v_w712_v);
	assign v_w5287_v = ~(v_w5286_v | v_w674_v);
	assign v_w2434_v = ~(v_w2399_v | v_w2318_v);
	assign v_w6059_v = ~(v_w6046_v | v_w6058_v);
	assign v_w2550_v = ~(v_w2150_v | v_w2287_v);
	assign v_w6566_v = ~(v_w6564_v & v_w6565_v);
	assign v_w6295_v = ~(v_w6293_v | v_w6294_v);
	assign v_w5072_v = ~(v_w5071_v & v_w673_v);
	assign v_w2612_v = ~(v_w8139_v);
	assign v_w4366_v = ~(v_w4362_v ^ v_w4365_v);
	assign v_w6539_v = ~(v_s400_v & v_w1701_v);
	assign v_w2946_v = ~(v_w2943_v | v_w2945_v);
	assign v_w3037_v = ~(v_s99_v & v_w565_v);
	assign v_w232_v = ~(v_w4056_v | v_w4082_v);
	assign v_w8251_v = v_w1008_v ^ v_w4577_v;
	assign v_w5284_v = ~(v_w2447_v & v_w3118_v);
	assign v_w254_v = ~(v_w5562_v & v_w5563_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s495_v<=0;
	end
	else
	begin
	v_s495_v<=v_w294_v;
	end
	end
	assign v_w6781_v = ~(v_s402_v & v_w656_v);
	assign v_w3528_v = ~(v_w3527_v);
	assign v_w178_v = ~(v_w5174_v & v_w5175_v);
	assign v_w3702_v = ~(v_w3700_v | v_w3701_v);
	assign v_w936_v = ~(v_w934_v | v_w935_v);
	assign v_w3646_v = ~(v_w3645_v);
	assign v_w6723_v = ~(v_w1734_v | v_w6579_v);
	assign v_w4378_v = ~(v_w4375_v | v_w4377_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s222_v<=0;
	end
	else
	begin
	v_s222_v<=v_w235_v;
	end
	end
	assign v_w6585_v = ~(v_w6583_v & v_w6584_v);
	assign v_w7016_v = v_w1592_v ^ v_w1028_v;
	assign v_w2547_v = ~(v_w2545_v | v_w2546_v);
	assign v_w163_v = v_s154_v & v_w5134_v;
	assign v_w2223_v = ~(v_s135_v | v_s134_v);
	assign v_w139_v = v_s130_v & v_w5134_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s79_v<=0;
	end
	else
	begin
	v_s79_v<=v_w87_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s247_v<=0;
	end
	else
	begin
	v_s247_v<=v_w260_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s472_v<=0;
	end
	else
	begin
	v_s472_v<=v_w525_v;
	end
	end
	assign v_w6036_v = ~(v_w6025_v & v_w6035_v);
	assign v_w6113_v = ~(v_w6111_v | v_w6112_v);
	assign v_w21_v = ~(v_w5614_v & v_w5615_v);
	assign v_w7687_v = ~(v_w831_v & v_w1783_v);
	assign v_w7749_v = ~(v_s121_v & v_w7742_v);
	assign v_w5212_v = ~(v_w693_v | v_w2883_v);
	assign v_w4213_v = ~(v_w2822_v ^ v_s210_v);
	assign v_w2227_v = ~(v_w2219_v & v_w2226_v);
	assign v_w884_v = ~(v_w882_v | v_w883_v);
	assign v_w1749_v = ~(v_w1297_v ^ v_w961_v);
	assign v_w784_v = ~(v_w8197_v);
	assign v_w6342_v = ~(v_s197_v & v_w6317_v);
	assign v_w7185_v = ~(v_w7183_v | v_w7184_v);
	assign v_w6930_v = ~(v_w1856_v | v_w6608_v);
	assign v_w7619_v = ~(v_w1739_v | v_w7618_v);
	assign v_w1713_v = ~(v_w1710_v | v_w1712_v);
	assign v_w488_v = ~(v_w5869_v & v_w5875_v);
	assign v_w7959_v = ~(v_s76_v & v_w2143_v);
	assign v_w4763_v = ~(v_w2448_v & v_w3025_v);
	assign v_w7221_v = ~(v_w7219_v | v_w7220_v);
	assign v_w4953_v = ~(v_w2914_v | v_w2370_v);
	assign v_w663_v = ~(v_w1972_v | v_w6012_v);
	assign v_w2895_v = ~(v_w1646_v | v_w2294_v);
	assign v_w1222_v = ~(v_w612_v & v_s393_v);
	assign v_w7995_v = ~(v_s464_v | v_s330_v);
	assign v_w2848_v = ~(v_w2847_v | v_w557_v);
	assign v_w5047_v = ~(v_w5040_v & v_w5046_v);
	assign v_w152_v = v_s143_v & v_w5134_v;
	assign v_w806_v = ~(v_w1109_v | v_w1059_v);
	assign v_w1151_v = v_s305_v | v_w1150_v;
	assign v_w7980_v = v_s472_v ^ v_s392_v;
	assign v_w1332_v = ~(v_w874_v & v_s414_v);
	assign v_w3301_v = ~(v_w3299_v & v_w3300_v);
	assign v_w4609_v = ~(v_w4608_v & v_w4582_v);
	assign v_w7286_v = ~(v_w7282_v & v_w7285_v);
	assign v_w6476_v = ~(v_w1407_v & v_w6019_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s487_v<=0;
	end
	else
	begin
	v_s487_v<=v_w175_v;
	end
	end
	assign v_w283_v = ~(v_w5094_v & v_w5095_v);
	assign v_w2454_v = ~(v_w2241_v & v_w865_v);
	assign v_w7998_v = ~(v_s462_v | v_s315_v);
	assign v_w5815_v = ~(v_w5809_v | v_w5814_v);
	assign v_w4845_v = ~(v_w2447_v & v_w2967_v);
	assign v_w4906_v = v_w4535_v ^ v_w4479_v;
	assign v_w7691_v = ~(v_w654_v & v_w7690_v);
	assign v_w1089_v = ~(v_w1420_v & v_w1426_v);
	assign v_w3216_v = ~(v_w2426_v);
	assign v_w1946_v = ~(v_w1944_v & v_w1945_v);
	assign v_w817_v = ~(v_w815_v | v_w816_v);
	assign v_w149_v = v_s140_v & v_w5134_v;
	assign v_w105_v = ~(v_w7784_v & v_w7785_v);
	assign v_w3908_v = v_w3902_v & v_w3905_v;
	assign v_w1300_v = ~(v_w1299_v & v_w809_v);
	assign v_w1675_v = ~(v_w1674_v | v_w1180_v);
	assign v_w7700_v = ~(v_w6995_v | v_w1919_v);
	assign v_w7692_v = ~(v_s235_v & v_w7667_v);
	assign v_w2923_v = ~(v_w697_v & v_w2922_v);
	assign v_w4303_v = ~(v_w4301_v & v_w4302_v);
	assign v_w4944_v = v_w2861_v ^ v_w4402_v;
	assign v_w3995_v = ~(v_w3994_v & v_w873_v);
	assign v_w5376_v = ~(v_w4954_v & v_w5375_v);
	assign v_w474_v = ~(v_w5668_v & v_w5669_v);
	assign v_w869_v = ~(v_w867_v | v_w868_v);
	assign v_w4765_v = ~(v_w4763_v & v_w4764_v);
	assign v_w6180_v = ~(v_w5977_v & v_w6179_v);
	assign v_w556_v = v_w8071_v ^ v_keyinput_7_v;
	assign v_w8157_v = v_w8156_v ^ v_keyinput_63_v;
	assign v_w7856_v = ~(v_s246_v & v_w1993_v);
	assign v_w6889_v = ~(v_w656_v & v_s344_v);
	assign v_w5684_v = ~(v_w613_v & v_s475_v);
	assign v_w4777_v = v_w4453_v ^ v_w4561_v;
	assign v_w1993_v = ~(v_w651_v);
	assign v_w2889_v = ~(v_w558_v & v_w1017_v);
	assign v_w6804_v = ~(v_w6803_v);
	assign v_w293_v = ~(v_w5254_v & v_w5255_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s435_v<=0;
	end
	else
	begin
	v_s435_v<=v_w487_v;
	end
	end
	assign v_w4519_v = ~(v_w871_v | v_w2671_v);
	assign v_w5958_v = ~(v_w2137_v & v_w578_v);
	assign v_w6122_v = ~(v_w6119_v | v_w6121_v);
	assign v_w3823_v = ~(v_w3521_v | v_w3735_v);
	assign v_w5398_v = ~(v_w5396_v & v_w5397_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s394_v<=0;
	end
	else
	begin
	v_s394_v<=v_w443_v;
	end
	end
	assign v_w5908_v = ~(v_w5904_v | v_w5907_v);
	assign v_w2086_v = v_w1324_v ^ v_w2000_v;
	assign v_w43_v = ~(v_w7915_v & v_w7916_v);
	assign v_w2653_v = v_w2652_v & v_s381_v;
	assign v_w685_v = v_s79_v ^ v_w1771_v;
	assign v_w4040_v = ~(v_w569_v | v_w4030_v);
	assign v_w6097_v = ~(v_w6074_v & v_w6073_v);
	assign v_w6937_v = ~(v_w6934_v | v_w6936_v);
	assign v_w3848_v = ~(v_w3846_v & v_w3847_v);
	assign v_w7066_v = ~(v_w596_v | v_w6579_v);
	assign v_w8000_v = ~(v_s460_v | v_s297_v);
	assign v_w7015_v = ~(v_w7013_v & v_w7014_v);
	assign v_w2575_v = ~(v_w2573_v & v_w2574_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s287_v<=0;
	end
	else
	begin
	v_s287_v<=v_w307_v;
	end
	end
	assign v_w7595_v = ~(v_w1762_v & v_w7245_v);
	assign v_w4856_v = ~(v_w2342_v | v_w4855_v);
	assign v_w984_v = ~(v_w2019_v | v_w1834_v);
	assign v_w7547_v = ~(v_w7258_v | v_w7546_v);
	assign v_w3295_v = ~(v_w3001_v ^ v_w3002_v);
	assign v_w415_v = ~(v_s512_v);
	assign v_w2257_v = ~(v_w2238_v & v_w879_v);
	assign v_w4459_v = ~(v_w3521_v & v_w2619_v);
	assign v_w4398_v = ~(v_w2296_v & v_w2339_v);
	assign v_w4718_v = ~(v_w674_v & v_s403_v);
	assign v_w4059_v = ~(v_w4057_v & v_w4058_v);
	assign v_w3222_v = ~(v_w2248_v & v_w3221_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s31_v<=0;
	end
	else
	begin
	v_s31_v<=v_w35_v;
	end
	end
	assign v_w7432_v = ~(v_w7387_v & v_w7431_v);
	assign v_w5258_v = ~(v_w5256_v | v_w5257_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s457_v<=0;
	end
	else
	begin
	v_s457_v<=v_w510_v;
	end
	end
	assign v_w5942_v = ~(v_w1343_v | v_w2135_v);
	assign v_w5448_v = ~(v_w4766_v | v_w5123_v);
	assign v_w520_v = ~(v_w6375_v & v_w6395_v);
	assign v_w2404_v = ~(v_w2402_v & v_w2403_v);
	assign v_w1326_v = ~(v_w1325_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s271_v<=0;
	end
	else
	begin
	v_s271_v<=v_w289_v;
	end
	end
	assign v_w1886_v = ~(v_w1884_v & v_w1885_v);
	assign v_w3184_v = ~(v_w3183_v & v_w3126_v);
	assign v_w2117_v = ~(v_w2115_v | v_w2116_v);
	assign v_w2077_v = ~(v_w2075_v | v_w2076_v);
	assign v_w3005_v = v_w425_v ^ v_w2650_v;
	assign v_w4222_v = ~(v_w2851_v | v_w4041_v);
	assign v_w173_v = ~(v_w5158_v & v_w5159_v);
	assign v_w687_v = v_w685_v & v_w686_v;
	assign v_w2196_v = ~(v_w2162_v);
	assign v_w3838_v = ~(v_w2368_v & v_w3731_v);
	assign v_w2733_v = ~(v_w2731_v & v_w2732_v);
	assign v_w3797_v = ~(v_w3794_v & v_w3796_v);
	assign v_w7624_v = ~(v_w7596_v & v_w7623_v);
	assign v_w5493_v = ~(v_w5491_v & v_w5492_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s158_v<=0;
	end
	else
	begin
	v_s158_v<=v_w167_v;
	end
	end
	assign v_w3755_v = ~(v_w753_v & v_w881_v);
	assign v_w271_v = ~(v_w5122_v & v_w5133_v);
	assign v_w4457_v = ~(v_w3638_v);
	assign v_w1207_v = ~(v_w1205_v & v_w1206_v);
	assign v_w3451_v = ~(v_w3449_v & v_w3450_v);
	assign v_w6578_v = ~(v_w1374_v & v_w1144_v);
	assign v_w4654_v = ~(v_w4653_v & v_w673_v);
	assign v_w3950_v = ~(v_w3940_v | v_w3949_v);
	assign v_w3127_v = ~(v_w3124_v & v_w3126_v);
	assign v_w6760_v = ~(v_w1718_v | v_w6571_v);
	assign v_w4318_v = ~(v_w2961_v & v_s118_v);
	assign v_w2071_v = ~(v_w2006_v | v_w2070_v);
	assign v_w7279_v = ~(v_w7275_v & v_w7278_v);
	assign v_w6021_v = ~(v_w6020_v);
	assign v_w1251_v = ~(v_w612_v & v_s318_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s241_v<=0;
	end
	else
	begin
	v_s241_v<=v_w254_v;
	end
	end
	assign v_w5438_v = ~(v_w5037_v & v_w4794_v);
	assign v_w6556_v = v_w6555_v ^ v_w6545_v;
	assign v_w6699_v = v_w1738_v ^ v_w1741_v;
	assign v_w4895_v = ~(v_w4893_v | v_w4894_v);
	assign v_w3225_v = ~(v_w3219_v | v_w3224_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s61_v<=0;
	end
	else
	begin
	v_s61_v<=v_w69_v;
	end
	end
	assign v_w7618_v = ~(v_w7597_v | v_w7617_v);
	assign v_w7782_v = ~(v_w7780_v | v_w7781_v);
	assign v_w5653_v = ~(v_w420_v & v_w2791_v);
	assign v_w3057_v = ~(v_w2361_v | v_w3056_v);
	assign v_w4513_v = ~(v_w4512_v & v_w3629_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s492_v<=0;
	end
	else
	begin
	v_s492_v<=v_w273_v;
	end
	end
	assign v_w4966_v = ~(v_w4965_v & v_w2456_v);
	assign v_w192_v = ~(v_w5426_v & v_w5433_v);
	assign v_w3220_v = ~(v_w2417_v & v_w2639_v);
	assign v_w1798_v = ~(v_w1797_v);
	assign v_w5621_v = ~(v_w420_v & v_w3216_v);
	assign v_w4780_v = ~(v_w4778_v & v_w4779_v);
	assign v_w3042_v = ~(v_w1078_v | v_w557_v);
	assign v_w920_v = ~(v_w919_v);
	assign v_w1965_v = ~(v_w1964_v | v_w8_v);
	assign v_w4540_v = ~(v_w3649_v & v_w4539_v);
	assign v_w5616_v = ~(v_s15_v & v_w676_v);
	assign v_w5230_v = ~(v_w5228_v | v_w5229_v);
	assign v_w270_v = ~(v_w5558_v & v_w5559_v);
	assign v_w5465_v = ~(v_w5463_v & v_w5464_v);
	assign v_w5651_v = ~(v_w420_v & v_w2993_v);
	assign v_w1778_v = ~(v_w1774_v | v_w1772_v);
	assign v_w5089_v = ~(v_w673_v & v_w5088_v);
	assign v_w7512_v = ~(v_w7504_v | v_w7511_v);
	assign v_w2458_v = ~(v_w674_v | v_w2457_v);
	assign v_w2524_v = ~(v_w2522_v | v_w2523_v);
	assign v_w620_v = v_w618_v & v_w619_v;
	assign v_w211_v = ~(v_w7937_v & v_w7938_v);
	assign v_w3798_v = ~(v_w3792_v & v_w3797_v);
	assign v_w2064_v = ~(v_w2063_v);
	assign v_w388_v = ~(v_w4905_v & v_w4915_v);
	assign v_w4325_v = ~(v_w2985_v & v_w887_v);
	assign v_w3895_v = ~(v_w3893_v & v_w3894_v);
	assign v_w1446_v = v_w373_v ^ v_w1157_v;
	assign v_w2959_v = ~(v_s476_v & v_w2778_v);
	assign v_w6086_v = ~(v_w6063_v | v_w6033_v);
	assign v_w4104_v = v_w4101_v ^ v_w4103_v;
	assign v_w4629_v = ~(v_w2448_v & v_w2690_v);
	assign v_w8085_v = v_w8084_v ^ v_keyinput_16_v;
	assign v_w4030_v = ~(v_w2193_v | v_w2242_v);
	assign v_w4604_v = ~(v_w3626_v ^ v_w4520_v);
	assign v_w7574_v = ~(v_w6802_v | v_w7573_v);
	assign v_w162_v = v_s153_v & v_w5134_v;
	assign v_w7896_v = ~(v_w651_v & v_w7795_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s184_v<=0;
	end
	else
	begin
	v_s184_v<=v_w197_v;
	end
	end
	assign v_w2769_v = ~(v_w2767_v & v_w2768_v);
	assign v_w5710_v = ~(v_w5708_v & v_w5709_v);
	assign v_w6244_v = ~(v_w6242_v & v_w6243_v);
	assign v_w1751_v = ~(v_w1286_v & v_w1003_v);
	assign v_w4727_v = ~(v_w4724_v | v_w4726_v);
	assign v_w5927_v = ~(v_w2009_v | v_w2010_v);
	assign v_w3281_v = ~(v_w3121_v | v_w2296_v);
	assign v_w7872_v = ~(v_s205_v & v_w1993_v);
	assign v_w4255_v = ~(v_w4253_v & v_w4254_v);
	assign v_w7104_v = ~(v_w7097_v & v_w7103_v);
	assign v_o15_v = ~(v_w8018_v ^ v_w8019_v);
	assign v_w5559_v = ~(v_w675_v & v_w5303_v);
	assign v_w7217_v = ~(v_w7215_v | v_w7216_v);
	assign v_w1964_v = ~(v_s79_v | v_w1771_v);
	assign v_w1911_v = v_w1909_v | v_w1910_v;
	assign v_w4761_v = v_w4563_v ^ v_w4452_v;
	assign v_w7966_v = ~(v_w527_v & v_w1309_v);
	assign v_w7267_v = ~(v_w687_v & v_w1309_v);
	assign v_w2111_v = ~(v_w2110_v & v_w2107_v);
	assign v_w276_v = ~(v_w3215_v & v_w3225_v);
	assign v_w3571_v = ~(v_w3566_v | v_w3570_v);
	assign v_w3930_v = ~(v_w3777_v & v_w3929_v);
	assign v_w3272_v = ~(v_w3270_v & v_w3271_v);
	assign v_w5601_v = ~(v_w5555_v & v_w5478_v);
	assign v_w1454_v = ~(v_w1445_v & v_w1453_v);
	assign v_w824_v = ~(v_w2294_v | v_w1664_v);
	assign v_w3169_v = ~(v_s277_v | v_w2635_v);
	assign v_w2904_v = ~(v_w699_v & v_s199_v);
	assign v_w2025_v = ~(v_w2018_v | v_w2024_v);
	assign v_w4241_v = ~(v_w2852_v & v_s202_v);
	assign v_w7142_v = ~(v_w7140_v | v_w7141_v);
	assign v_w7197_v = ~(v_w7195_v | v_w7196_v);
	assign v_w4026_v = ~(v_w4025_v & v_w554_v);
	assign v_w969_v = ~(v_in19_v ^ v_w1235_v);
	assign v_w4484_v = ~(v_w2890_v | v_w1017_v);
	assign v_w7077_v = ~(v_w7075_v & v_w7076_v);
	assign v_w3573_v = ~(v_w2706_v | v_w754_v);
	assign v_w3751_v = v_w3595_v & v_w881_v;
	assign v_w1819_v = ~(v_w901_v & v_w1445_v);
	assign v_w842_v = ~(v_w840_v | v_w841_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s368_v<=0;
	end
	else
	begin
	v_s368_v<=v_w411_v;
	end
	end
	assign v_w2157_v = v_w2156_v & v_s476_v;
	assign v_w6329_v = ~(v_s324_v & v_w1626_v);
	assign v_w1608_v = ~(v_s318_v & v_w562_v);
	assign v_w811_v = ~(v_w2693_v ^ v_w2696_v);
	assign v_w5711_v = ~(v_w5706_v | v_w5710_v);
	assign v_w4052_v = ~(v_w4047_v | v_w4051_v);
	assign v_w1830_v = ~(v_w578_v);
	assign v_w2104_v = ~(v_w2101_v ^ v_w2103_v);
	assign v_w4887_v = ~(v_w4884_v | v_w4886_v);
	assign v_w7330_v = ~(v_w679_v | v_w1091_v);
	assign v_w8224_v = v_w8223_v ^ v_keyinput_109_v;
	assign v_w58_v = v_s50_v & v_w7107_v;
	assign v_w517_v = ~(v_w6292_v & v_w6313_v);
	assign v_w2795_v = ~(v_w1476_v | v_w2294_v);
	assign v_w333_v = ~(v_w5238_v & v_w5239_v);
	assign v_w6709_v = ~(v_w1798_v & v_w1337_v);
	assign v_w5536_v = ~(v_w5276_v & v_w5126_v);
	assign v_w5246_v = ~(v_w5244_v | v_w5245_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s490_v<=0;
	end
	else
	begin
	v_s490_v<=v_w262_v;
	end
	end
	assign v_w7552_v = ~(v_w7550_v | v_w7551_v);
	assign v_w2844_v = ~(v_w2358_v & v_s329_v);
	assign v_w8083_v = v_w8082_v ^ v_keyinput_15_v;
	assign v_w6783_v = ~(v_w1140_v & v_w1696_v);
	assign v_w1844_v = ~(v_w1831_v & v_w1843_v);
	assign v_w2123_v = ~(v_w2122_v);
	assign v_w2913_v = v_w552_v ^ v_w2912_v;
	assign v_w2396_v = ~(v_s277_v | v_w2361_v);
	assign v_w1283_v = ~(v_w1052_v & v_s447_v);
	assign v_w7950_v = ~(v_w527_v & v_w1401_v);
	assign v_w7779_v = ~(v_s101_v & v_w7742_v);
	assign v_w6365_v = ~(v_w5808_v & v_w6364_v);
	assign v_w7912_v = ~(v_w651_v & v_w7845_v);
	assign v_w2098_v = ~(v_w8135_v);
	assign v_w2116_v = ~(v_w1918_v | v_w2109_v);
	assign v_w5346_v = ~(v_w683_v & v_w5345_v);
	assign v_w7161_v = ~(v_w7159_v | v_w7160_v);
	assign v_w4536_v = v_w2382_v & v_w2444_v;
	assign v_w700_v = ~(v_w2165_v | v_w2176_v);
	assign v_w6913_v = ~(v_w6911_v & v_w6912_v);
	assign v_w593_v = ~(v_w544_v | v_w592_v);
	assign v_w1490_v = ~(v_s301_v ^ v_w1489_v);
	assign v_w5596_v = ~(v_s94_v & v_w676_v);
	assign v_w1256_v = ~(v_s309_v & v_w1192_v);
	assign v_w505_v = ~(v_w6588_v & v_w6589_v);
	assign v_w5005_v = ~(v_w4994_v | v_w5004_v);
	assign v_w4031_v = ~(v_w2235_v & v_w4030_v);
	assign v_w2105_v = ~(v_w1963_v | v_w1981_v);
	assign v_w6643_v = ~(v_w6641_v & v_w6642_v);
	assign v_w1590_v = ~(v_w1588_v | v_w1589_v);
	assign v_w7586_v = ~(v_w2102_v | v_w7585_v);
	assign v_w6044_v = ~(v_w664_v & v_s455_v);
	assign v_w3458_v = ~(v_w612_v & v_s16_v);
	assign v_w4188_v = ~(v_w4173_v & v_w4176_v);
	assign v_w7770_v = ~(v_w7768_v | v_w7769_v);
	assign v_w1926_v = ~(v_w1925_v);
	assign v_w4427_v = ~(v_w3468_v | v_w2264_v);
	assign v_w7873_v = ~(v_w651_v & v_w7728_v);
	assign v_w3231_v = ~(v_w621_v | v_w2729_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s7_v<=0;
	end
	else
	begin
	v_s7_v<=v_w7_v;
	end
	end
	assign v_w2563_v = ~(v_w2562_v | v_w617_v);
	assign v_w458_v = ~(v_w6742_v & v_w6743_v);
	assign v_w3942_v = ~(v_w3936_v | v_w1011_v);
	assign v_w7018_v = ~(v_w7015_v | v_w7017_v);
	assign v_w622_v = ~(v_w2729_v | v_w3051_v);
	assign v_w7521_v = ~(v_w7272_v & v_w7520_v);
	assign v_w5009_v = ~(v_w2265_v & v_w2575_v);
	assign v_w8180_v = v_w8179_v ^ v_keyinput_82_v;
	assign v_w7461_v = ~(v_w1624_v | v_w680_v);
	assign v_w4203_v = v_w4199_v ^ v_w4202_v;
	assign v_w1670_v = ~(v_w562_v & v_s120_v);
	assign v_w1096_v = ~(v_w1095_v);
	assign v_w904_v = ~(v_w2041_v & v_w2045_v);
	assign v_w56_v = v_s48_v & v_w7107_v;
	assign v_w4998_v = v_w4539_v ^ v_w3649_v;
	assign v_w8232_v = v_w8231_v ^ v_keyinput_115_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s208_v<=0;
	end
	else
	begin
	v_s208_v<=v_w221_v;
	end
	end
	assign v_w2681_v = ~(v_w2676_v | v_w2680_v);
	assign v_w2474_v = ~(v_w2472_v | v_w2473_v);
	assign v_w2830_v = v_w552_v ^ v_w2829_v;
	assign v_w5114_v = ~(v_w2331_v | v_w2264_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s106_v<=0;
	end
	else
	begin
	v_s106_v<=v_w114_v;
	end
	end
	assign v_w3637_v = ~(v_w3559_v & v_w3565_v);
	assign v_w598_v = v_w600_v & v_w601_v;
	assign v_w4259_v = ~(v_w2929_v ^ v_s350_v);
	assign v_w5788_v = ~(v_w892_v & v_w1835_v);
	assign v_w3974_v = ~(v_w3972_v & v_w3973_v);
	assign v_w4667_v = ~(v_w4665_v & v_w4666_v);
	assign v_w1905_v = ~(v_w1297_v & v_w961_v);
	assign v_w1059_v = ~(v_w842_v | v_w1058_v);
	assign v_w4339_v = ~(v_s117_v & v_w4320_v);
	assign v_w5341_v = ~(v_w4863_v | v_w5031_v);
	assign v_w5315_v = ~(v_w5054_v & v_w5037_v);
	assign v_w7925_v = ~(v_s289_v & v_w6015_v);
	assign v_w696_v = ~(v_w2354_v & v_w544_v);
	assign v_w8048_v = ~(v_w7982_v | v_w8047_v);
	assign v_w2328_v = ~(v_w563_v & v_s87_v);
	assign v_w1609_v = ~(v_w715_v | v_w8_v);
	assign v_w4206_v = ~(v_w3323_v & v_w4205_v);
	assign v_w4608_v = ~(v_w4607_v & v_w3626_v);
	assign v_w3261_v = ~(v_w3258_v & v_w3260_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s14_v<=0;
	end
	else
	begin
	v_s14_v<=v_w15_v;
	end
	end
	assign v_w5173_v = v_w5141_v & v_s38_v;
	assign v_w434_v = ~(v_w3428_v & v_w3435_v);
	assign v_w4082_v = ~(v_w695_v);
	assign v_w5606_v = ~(v_s39_v & v_w676_v);
	assign v_w6359_v = ~(v_s338_v & v_w6332_v);
	assign v_w5403_v = ~(v_s176_v & v_w5386_v);
	assign v_w2409_v = ~(v_w2407_v & v_w2408_v);
	assign v_w6383_v = ~(v_w6029_v | v_w6382_v);
	assign v_w7009_v = ~(v_w6592_v & v_w789_v);
	assign v_w1790_v = ~(v_w759_v & v_w1789_v);
	assign v_w3499_v = ~(v_w3498_v | v_w2418_v);
	assign v_w6075_v = ~(v_w6073_v ^ v_w6074_v);
	assign v_w6998_v = ~(v_w1848_v ^ v_w790_v);
	assign v_w3828_v = v_w3826_v | v_w3827_v;
	assign v_w8065_v = ~(v_w3041_v | v_w3044_v);
	assign v_w8138_v = ~(v_w2610_v & v_w2611_v);
	assign v_w4210_v = ~(v_w4208_v & v_w4209_v);
	assign v_w5907_v = ~(v_w5906_v | v_w5693_v);
	assign v_w1377_v = ~(v_w1376_v | v_w8_v);
	assign v_w7041_v = ~(v_w7039_v & v_w7040_v);
	assign v_w1999_v = v_w723_v;
	assign v_w703_v = ~(v_w546_v & v_w785_v);
	assign v_w3257_v = ~(v_w3255_v | v_w3256_v);
	assign v_w6163_v = ~(v_w6162_v & v_w659_v);
	assign v_w5062_v = ~(v_w8161_v);
	assign v_w4179_v = ~(v_w4172_v & v_w4178_v);
	assign v_w5317_v = ~(v_w5315_v & v_w5316_v);
	assign v_w3123_v = ~(v_w3120_v | v_w3122_v);
	assign v_w4069_v = ~(v_w690_v & v_w4068_v);
	assign v_w823_v = ~(v_w2876_v & v_w2885_v);
	assign v_w5795_v = ~(v_w5793_v & v_w5794_v);
	assign v_w5929_v = ~(v_w5928_v & v_w2113_v);
	assign v_w1217_v = ~(v_w1215_v & v_w1216_v);
	assign v_w6270_v = ~(v_w657_v & v_s322_v);
	assign v_w5898_v = ~(v_w5895_v ^ v_w5897_v);
	assign v_w4218_v = ~(v_w4217_v & v_w692_v);
	assign v_w137_v = v_s128_v & v_w5134_v;
	assign v_w6784_v = ~(v_w6782_v & v_w6783_v);
	assign v_w3101_v = ~(v_w558_v & v_w3100_v);
	assign v_w5625_v = ~(v_w420_v & v_w1131_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s399_v<=0;
	end
	else
	begin
	v_s399_v<=v_w448_v;
	end
	end
	assign v_w6202_v = ~(v_w6172_v & v_w6201_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s507_v<=0;
	end
	else
	begin
	v_s507_v<=v_w383_v;
	end
	end
	assign v_w133_v = ~(v_w5214_v & v_w5215_v);
	assign v_w1616_v = v_w8158_v ^ v_keyinput_64_v;
	assign v_w603_v = ~(v_w602_v ^ v_w596_v);
	assign v_w4352_v = ~(v_w3289_v & v_w4351_v);
	assign v_w2399_v = ~(v_w2397_v & v_w2398_v);
	assign v_w7919_v = ~(v_s248_v & v_w6015_v);
	assign v_w5899_v = ~(v_w5693_v | v_w5898_v);
	assign v_w3322_v = ~(v_w3320_v | v_w3321_v);
	assign v_w88_v = ~(v_w7796_v & v_w7797_v);
	assign v_w7611_v = ~(v_w7609_v | v_w7610_v);
	assign v_w4006_v = v_w8181_v ^ v_keyinput_83_v;
	assign v_w2150_v = ~(v_s290_v | v_s291_v);
	assign v_w431_v = ~(v_w3307_v & v_w3308_v);
	assign v_w4346_v = ~(v_w2756_v ^ v_s106_v);
	assign v_w4595_v = ~(v_w2660_v & v_w2347_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s420_v<=0;
	end
	else
	begin
	v_s420_v<=v_w471_v;
	end
	end
	assign v_w2760_v = v_w552_v ^ v_w2759_v;
	assign v_w6080_v = ~(v_w6078_v & v_w6079_v);
	assign v_w6667_v = ~(v_w1787_v & v_w1323_v);
	assign v_w5610_v = ~(v_s28_v & v_w676_v);
	assign v_w7118_v = ~(v_w7117_v);
	assign v_w2500_v = ~(v_w2498_v & v_w2499_v);
	assign v_w7813_v = ~(v_w7811_v | v_w7812_v);
	assign v_w1320_v = ~(v_w1318_v & v_w1319_v);
	assign v_w625_v = ~(v_w623_v | v_w624_v);
	assign v_w1606_v = ~(v_w1604_v & v_w1605_v);
	assign v_w816_v = ~(v_w3082_v & v_w3083_v);
	assign v_w6927_v = ~(v_w6925_v & v_w6926_v);
	assign v_w1991_v = ~(v_w1990_v & v_w1987_v);
	assign v_w4681_v = ~(v_w4680_v & v_w878_v);
	assign v_w3389_v = ~(v_w3387_v & v_w3388_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s141_v<=0;
	end
	else
	begin
	v_s141_v<=v_w150_v;
	end
	end
	assign v_w369_v = ~(v_w6921_v & v_w6928_v);
	assign v_w1427_v = ~(v_w736_v ^ v_w1272_v);
	assign v_w1178_v = ~(v_w780_v | v_s424_v);
	assign v_w5466_v = ~(v_w4725_v | v_w5123_v);
	assign v_w4957_v = v_s316_v & v_w674_v;
	assign v_w2762_v = ~(v_w2484_v & v_w2761_v);
	assign v_w2692_v = ~(v_w2682_v & v_w2691_v);
	assign v_w4343_v = ~(v_w4337_v | v_w4340_v);
	assign v_w1657_v = ~(v_w1655_v | v_w1656_v);
	assign v_w3485_v = ~(v_w3199_v);
	assign v_w1040_v = ~(v_s36_v & v_w1104_v);
	assign v_w8141_v = v_w8140_v ^ v_keyinput_52_v;
	assign v_w348_v = ~(v_w6946_v & v_w6961_v);
	assign v_w3382_v = v_w8090_v ^ v_keyinput_19_v;
	assign v_w2767_v = ~(v_w8200_v);
	assign v_w1142_v = v_w1103_v & v_s6_v;
	assign v_w127_v = ~(v_w5584_v & v_w5585_v);
	assign v_w309_v = ~(v_w7925_v & v_w7926_v);
	assign v_w7058_v = ~(v_w7056_v | v_w7057_v);
	assign v_w375_v = ~(v_w6003_v & v_w6010_v);
	assign v_w4864_v = ~(v_w2965_v ^ v_w4406_v);
	assign v_w6926_v = ~(v_w1798_v & v_w1126_v);
	assign v_w7403_v = ~(v_w7398_v & v_w7401_v);
	assign v_w4790_v = ~(v_w4788_v | v_w4789_v);
	assign v_w6239_v = ~(v_w6237_v ^ v_w6238_v);
	assign v_w1508_v = ~(v_w1507_v | v_w1180_v);
	assign v_w2996_v = ~(v_w2972_v ^ v_w2989_v);
	assign v_w4521_v = ~(v_w3627_v | v_w4520_v);
	assign v_w6490_v = v_w1391_v ^ v_w6489_v;
	assign v_w3683_v = ~(v_w3624_v | v_w3682_v);
	assign v_w6146_v = v_w8093_v ^ v_keyinput_21_v;
	assign v_w326_v = ~(v_w5983_v & v_w5987_v);
	assign v_w4492_v = ~(v_w4456_v | v_w4491_v);
	assign v_w228_v = ~(v_w7868_v & v_w7869_v);
	assign v_w7311_v = ~(v_w680_v | v_w1074_v);
	assign v_w7549_v = ~(v_w7547_v | v_w7548_v);
	assign v_w4420_v = ~(v_w3087_v & v_w4419_v);
	assign v_w6407_v = v_w6399_v & v_w6405_v;
	assign v_w310_v = ~(v_w5246_v & v_w5247_v);
	assign v_w7121_v = ~(v_w528_v | v_w730_v);
	assign v_w6911_v = ~(v_w1612_v | v_w6910_v);
	assign v_w5074_v = ~(v_w5058_v | v_w5073_v);
	assign v_w6632_v = ~(v_w6630_v & v_w6631_v);
	assign v_w6618_v = ~(v_w6616_v & v_w6617_v);
	assign v_w944_v = ~(v_w1534_v & v_w1535_v);
	assign v_w3251_v = ~(v_w3121_v | v_w572_v);
	assign v_w2604_v = ~(v_s293_v & v_w693_v);
	assign v_w2118_v = ~(v_w1966_v | v_w528_v);
	assign v_w4881_v = ~(v_w825_v | v_w2264_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s259_v<=0;
	end
	else
	begin
	v_s259_v<=v_w275_v;
	end
	end
	assign v_w988_v = ~(v_w1506_v | v_w808_v);
	assign v_w1381_v = ~(v_w808_v | v_w1380_v);
	assign v_w4798_v = ~(v_w3012_v | v_w2370_v);
	assign v_w5443_v = ~(v_w683_v & v_w5442_v);
	assign v_w3682_v = ~(v_w3625_v & v_w3681_v);
	assign v_w5537_v = ~(v_w5535_v & v_w5536_v);
	assign v_w7034_v = ~(v_w7032_v | v_w7033_v);
	assign v_w6052_v = ~(v_w6051_v & v_w659_v);
	assign v_w4025_v = ~(v_w3730_v & v_w4024_v);
	assign v_w6233_v = ~(v_w664_v & v_s462_v);
	assign v_w3714_v = ~(v_w3713_v & v_w3565_v);
	assign v_w6928_v = ~(v_w655_v & v_w6927_v);
	assign v_w6931_v = ~(v_w6929_v | v_w6930_v);
	assign v_w7953_v = ~(v_s99_v & v_w2143_v);
	assign v_w7294_v = ~(v_w7286_v & v_w7293_v);
	assign v_w5737_v = ~(v_w5735_v | v_w5736_v);
	assign v_w6521_v = ~(v_s109_v & v_w6484_v);
	assign v_w5412_v = ~(v_w1083_v | v_w2602_v);
	assign v_w5104_v = v_w2427_v ^ v_w2461_v;
	assign v_w8131_v = v_w8130_v ^ v_keyinput_47_v;
	assign v_w1692_v = ~(v_w1052_v & v_s102_v);
	assign v_w1862_v = ~(v_w1860_v | v_w1861_v);
	assign v_w4830_v = ~(v_w4822_v | v_w4589_v);
	assign v_w3981_v = ~(v_w3979_v | v_w3980_v);
	assign v_w2302_v = ~(v_w565_v & v_s237_v);
	assign v_w1931_v = ~(v_w1930_v ^ v_s432_v);
	assign v_w7135_v = ~(v_w7118_v & v_w1289_v);
	assign v_w7316_v = ~(v_w7314_v | v_w7315_v);
	assign v_w2315_v = ~(v_w2310_v | v_w2314_v);
	assign v_w3287_v = ~(v_w3012_v | v_w2620_v);
	assign v_w4436_v = ~(v_w4434_v & v_w4435_v);
	assign v_w7808_v = ~(v_w654_v & v_w7807_v);
	assign v_w5880_v = ~(v_w2117_v & v_w831_v);
	assign v_w2813_v = ~(v_w2358_v & v_s316_v);
	assign v_w3698_v = ~(v_w3515_v | v_w3697_v);
	assign v_w7888_v = ~(v_w651_v & v_w7771_v);
	assign v_w4347_v = ~(v_s116_v & v_w2784_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s23_v<=0;
	end
	else
	begin
	v_s23_v<=v_w25_v;
	end
	end
	assign v_w1246_v = ~(v_s325_v & v_w1103_v);
	assign v_w6609_v = ~(v_w6601_v & v_w1114_v);
	assign v_w4551_v = ~(v_w3491_v | v_w4550_v);
	assign v_w3338_v = ~(v_w3035_v);
	assign v_w3665_v = ~(v_w3554_v & v_w3664_v);
	assign v_w5564_v = ~(v_s239_v & v_w676_v);
	assign v_w6983_v = v_w980_v ^ v_w1850_v;
	assign v_w5440_v = ~(v_w4781_v | v_w5123_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s104_v<=0;
	end
	else
	begin
	v_s104_v<=v_w112_v;
	end
	end
	assign v_w2087_v = ~(v_w2085_v | v_w2086_v);
	assign v_w6330_v = ~(v_w6290_v & v_w6289_v);
	assign v_w765_v = ~(v_w835_v | v_w836_v);
	assign v_w923_v = ~(v_w921_v | v_w922_v);
	assign v_w7177_v = ~(v_w7175_v | v_w7176_v);
	assign v_w3706_v = ~(v_w3704_v | v_w3705_v);
	assign v_w2175_v = v_w2174_v | v_s218_v;
	assign v_w6509_v = ~(v_w657_v & v_s400_v);
	assign v_w4768_v = ~(v_w4765_v | v_w4767_v);
	assign v_w1227_v = ~(v_s90_v & v_w1192_v);
	assign v_w5053_v = ~(v_w5051_v | v_w5052_v);
	assign v_w3678_v = ~(v_w3610_v | v_w3488_v);
	assign v_w159_v = v_s150_v & v_w5134_v;
	assign v_w7093_v = ~(v_w1140_v & v_s247_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s248_v<=0;
	end
	else
	begin
	v_s248_v<=v_w261_v;
	end
	end
	assign v_w1643_v = ~(v_w718_v | v_w8_v);
	assign v_w217_v = ~(v_w7729_v & v_w7730_v);
	assign v_w6218_v = v_w1490_v ^ v_w6217_v;
	assign v_w7275_v = ~(v_w7273_v & v_w7274_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s246_v<=0;
	end
	else
	begin
	v_s246_v<=v_w259_v;
	end
	end
	assign v_w3487_v = ~(v_w2300_v & v_w1767_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s69_v<=0;
	end
	else
	begin
	v_s69_v<=v_w77_v;
	end
	end
	assign v_w7858_v = ~(v_s244_v & v_w1993_v);
	assign v_w6831_v = ~(v_w6828_v & v_w6830_v);
	assign v_w3391_v = ~(v_w3389_v | v_w3390_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s503_v<=0;
	end
	else
	begin
	v_s503_v<=v_w364_v;
	end
	end
	assign v_w2716_v = ~(v_w2358_v & v_s403_v);
	assign v_w6403_v = ~(v_s160_v & v_w888_v);
	assign v_w5759_v = ~(v_w5757_v | v_w5758_v);
	assign v_w5518_v = ~(v_w3087_v | v_w2602_v);
	assign v_w2747_v = ~(v_w2358_v & v_s389_v);
	assign v_w3358_v = ~(v_w3357_v & v_w2947_v);
	assign v_w7506_v = ~(v_w680_v | v_w917_v);
	assign v_w5121_v = ~(v_w2335_v | v_w5120_v);
	assign v_w2016_v = ~(v_w596_v);
	assign v_w6812_v = ~(v_w1787_v & v_w1416_v);
	assign v_w5800_v = ~(v_w5799_v & v_w2113_v);
	assign v_w8005_v = ~(v_s377_v & v_s456_v);
	assign v_w606_v = ~(v_w1562_v | v_w1564_v);
	assign v_w5966_v = ~(v_w1816_v | v_w5734_v);
	assign v_w1415_v = ~(v_w1052_v & v_s89_v);
	assign v_w5260_v = ~(v_w1_v | v_w2330_v);
	assign v_w5889_v = ~(v_w2137_v & v_w1824_v);
	assign v_w2156_v = ~(v_w2146_v & v_w707_v);
	assign v_w4442_v = ~(v_w964_v | v_w2264_v);
	assign v_w1273_v = v_in15_v ^ v_w1223_v;
	assign v_w3080_v = v_w553_v ^ v_w3079_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s265_v<=0;
	end
	else
	begin
	v_s265_v<=v_w282_v;
	end
	end
	assign v_w4501_v = ~(v_w3338_v | v_w3177_v);
	assign v_w7793_v = ~(v_w6738_v | v_w7792_v);
	assign v_w6640_v = ~(v_w6639_v);
	assign v_w7891_v = ~(v_s98_v & v_w7876_v);
	assign v_w3277_v = ~(v_w3275_v & v_w3276_v);
	assign v_w952_v = ~(v_w920_v & v_w1135_v);
	assign v_w2381_v = ~(v_w2378_v | v_w2297_v);
	assign v_w4399_v = ~(v_w2558_v | v_w4398_v);
	assign v_w6891_v = ~(v_w6889_v & v_w6890_v);
	assign v_w4284_v = ~(v_w4275_v | v_w4283_v);
	assign v_w6223_v = ~(v_s224_v & v_w889_v);
	assign v_w3633_v = ~(v_w3578_v & v_w3569_v);
	assign v_w7865_v = ~(v_w651_v & v_w7703_v);
	assign v_w2414_v = ~(v_s255_v & v_w593_v);
	assign v_w5887_v = ~(v_w5885_v | v_w5886_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s286_v<=0;
	end
	else
	begin
	v_s286_v<=v_w306_v;
	end
	end
	assign v_w1553_v = ~(v_s270_v & v_w870_v);
	assign v_w4739_v = ~(v_w761_v | v_w2264_v);
	assign v_w3636_v = ~(v_w8229_v);
	assign v_w7939_v = ~(v_s346_v & v_w2143_v);
	assign v_w5374_v = ~(v_w5372_v & v_w5373_v);
	assign v_w1367_v = ~(v_s401_v ^ v_w1162_v);
	assign v_w6285_v = ~(v_w6280_v & v_w6284_v);
	assign v_w7659_v = ~(v_w7657_v & v_w7658_v);
	assign v_w2643_v = ~(v_w2642_v | v_w355_v);
	assign v_w3130_v = ~(v_w3109_v & v_w2993_v);
	assign v_w7368_v = ~(v_w7366_v | v_w7367_v);
	assign v_w4842_v = ~(v_w4840_v | v_w4841_v);
	assign v_w6249_v = ~(v_w1490_v & v_w6225_v);
	assign v_w2866_v = ~(v_w2860_v | v_w2865_v);
	assign v_w2437_v = ~(v_w2433_v | v_w2436_v);
	assign v_w7927_v = ~(v_s227_v & v_w6015_v);
	assign v_w7800_v = ~(v_w7798_v | v_w7799_v);
	assign v_w8024_v = ~(v_w8000_v | v_w8023_v);
	assign v_w2052_v = ~(v_w1650_v ^ v_w1999_v);
	assign v_w5857_v = ~(v_w597_v | v_w2062_v);
	assign v_w3079_v = ~(v_w3069_v & v_w3078_v);
	assign v_w4938_v = ~(v_w4936_v | v_w4937_v);
	assign v_w971_v = v_w970_v & v_w902_v;
	assign v_w2037_v = ~(v_w8224_v);
	assign v_w3454_v = ~(v_s4_v & v_w1192_v);
	assign v_w8150_v = ~(v_w4356_v ^ v_w4357_v);
	assign v_w3687_v = ~(v_w3686_v & v_w3480_v);
	assign v_w8201_v = v_w6660_v ^ v_keyinput_96_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s258_v<=0;
	end
	else
	begin
	v_s258_v<=v_w273_v;
	end
	end
	assign v_w1593_v = ~(v_w1592_v | v_w1028_v);
	assign v_w8118_v = v_w8117_v ^ v_keyinput_39_v;
	assign v_w6184_v = v_s304_v ^ v_w1503_v;
	assign v_w4070_v = ~(v_w887_v & v_w2321_v);
	assign v_w5558_v = ~(v_s255_v & v_w676_v);
	assign v_w1144_v = v_w1142_v | v_w1143_v;
	assign v_w6906_v = ~(v_w656_v & v_s338_v);
	assign v_w4602_v = ~(v_w2369_v & v_w3118_v);
	assign v_w7735_v = ~(v_w654_v & v_w7734_v);
	assign v_w7249_v = ~(v_w7244_v & v_w7248_v);
	assign v_w6363_v = ~(v_w6362_v & v_w6020_v);
	assign v_w6390_v = ~(v_w664_v & v_s467_v);
	assign v_w615_v = ~(v_w612_v | v_w613_v);
	assign v_w4289_v = v_w4285_v ^ v_w4288_v;
	assign v_w7943_v = ~(v_s161_v & v_w2143_v);
	assign v_w7748_v = ~(v_w654_v & v_w7747_v);
	assign v_w480_v = ~(v_w4530_v & v_w4593_v);
	assign v_w7012_v = ~(v_w7010_v | v_w7011_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s253_v<=0;
	end
	else
	begin
	v_s253_v<=v_w268_v;
	end
	end
	assign v_w1189_v = ~(v_w717_v | v_w8_v);
	assign v_w2939_v = v_w2936_v & v_w2938_v;
	assign v_w710_v = ~(v_w548_v | v_w560_v);
	assign v_w4542_v = ~(v_w3644_v & v_w4541_v);
	assign v_w734_v = ~(v_in19_v | v_w1235_v);
	assign v_w7083_v = ~(v_w6602_v | v_w7082_v);
	assign v_w7592_v = v_w7591_v ^ v_w1378_v;
	assign v_w8115_v = ~(v_w5252_v | v_w5253_v);
	assign v_w5020_v = ~(v_w3648_v | v_w4537_v);
	assign v_w8165_v = v_w3585_v & v_w3716_v;
	assign v_w7054_v = ~(v_w7050_v | v_w7053_v);
	assign v_w3245_v = ~(v_w636_v & v_w3244_v);
	assign v_w1705_v = ~(v_w1702_v | v_w1704_v);
	assign v_w5560_v = ~(v_s253_v & v_w676_v);
	assign v_w2859_v = v_w552_v ^ v_w2858_v;
	assign v_w7725_v = ~(v_w7693_v | v_w6935_v);
	assign v_w29_v = ~(v_w7903_v & v_w7904_v);
	assign v_w2332_v = ~(v_s36_v ^ v_w1104_v);
	assign v_w5357_v = ~(v_w4983_v | v_w5356_v);
	assign v_w8155_v = v_w8154_v ^ v_keyinput_62_v;
	assign v_w6530_v = v_w6526_v ^ v_w6529_v;
	assign v_w2254_v = ~(v_s167_v | v_w2199_v);
	assign v_w4499_v = ~(v_w4497_v | v_w4498_v);
	assign v_w1465_v = ~(v_s336_v ^ v_w1464_v);
	assign v_w3342_v = ~(v_w2722_v);
	assign v_w7850_v = ~(v_w654_v & v_w7849_v);
	assign v_w2717_v = ~(v_w2715_v & v_w2716_v);
	assign v_w3045_v = ~(v_w3041_v & v_w3044_v);
	assign v_w5078_v = ~(v_w2263_v & v_w2327_v);
	assign v_w3076_v = ~(v_w593_v & v_s42_v);
	assign v_w6557_v = ~(v_w6556_v & v_w659_v);
	assign v_w2400_v = ~(v_w2399_v);
	assign v_w6701_v = ~(v_w6698_v | v_w6700_v);
	assign v_w3016_v = ~(v_w3015_v | v_w531_v);
	assign v_w8214_v = v_w8213_v ^ v_keyinput_104_v;
	assign v_w6131_v = v_s236_v ^ v_w1528_v;
	assign v_w4105_v = ~(v_w4104_v & v_w692_v);
	assign v_w3590_v = ~(v_w3588_v | v_w3589_v);
	assign v_w3297_v = ~(v_w2635_v | v_w2702_v);
	assign v_w6642_v = v_w1748_v ^ v_w1749_v;
	assign v_w4972_v = ~(v_w4970_v | v_w4971_v);
	assign v_w5268_v = ~(v_w5266_v & v_w5267_v);
	assign v_w658_v = ~(v_w6013_v);
	assign v_w2229_v = ~(v_w2207_v & v_w2228_v);
	assign v_w4435_v = ~(v_w674_v & v_s426_v);
	assign v_w2503_v = ~(v_w2501_v | v_w2502_v);
	assign v_w439_v = ~(v_w4350_v & v_w4361_v);
	assign v_w2932_v = ~(v_w572_v | v_w617_v);
	assign v_w4429_v = ~(v_w1136_v & v_s40_v);
	assign v_w4925_v = ~(v_w4923_v & v_w4924_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s389_v<=0;
	end
	else
	begin
	v_s389_v<=v_w438_v;
	end
	end
	assign v_w2240_v = ~(v_w2239_v & v_s476_v);
	assign v_w4432_v = ~(v_w4431_v & v_w673_v);
	assign v_w3614_v = ~(v_w3609_v & v_w3613_v);
	assign v_w6670_v = ~(v_w6666_v | v_w6669_v);
	assign v_w2857_v = ~(v_w2856_v | v_w617_v);
	assign v_w4580_v = ~(v_w1006_v | v_w4579_v);
	assign v_w4933_v = v_w2901_v ^ v_w4403_v;
	assign v_w6398_v = ~(v_w6396_v & v_w6397_v);
	assign v_w1047_v = ~(v_w1044_v & v_w1273_v);
	assign v_w2689_v = ~(v_w699_v & v_s186_v);
	assign v_w7660_v = ~(v_w6638_v & v_w1919_v);
	assign v_w7241_v = ~(v_w7239_v & v_w7240_v);
	assign v_w7179_v = ~(v_w6399_v | v_w529_v);
	assign v_w6307_v = ~(v_w6306_v & v_w659_v);
	assign v_w1554_v = ~(v_w1552_v & v_w1553_v);
	assign v_w7964_v = ~(v_w527_v & v_w1323_v);
	assign v_w4899_v = ~(v_w572_v | v_w2264_v);
	assign v_w626_v = ~(v_w971_v & v_w2059_v);
	assign v_w4410_v = ~(v_w1011_v & v_w4409_v);
	assign v_w1061_v = ~(v_w805_v | v_w1060_v);
	assign v_w5257_v = ~(v_w2322_v | v_w1_v);
	assign v_w535_v = ~(v_w1582_v | v_w808_v);
	assign v_w3365_v = ~(v_w3363_v | v_w3364_v);
	assign v_w7920_v = ~(v_w527_v & v_w602_v);
	assign v_w142_v = v_s133_v & v_w5134_v;
	assign v_w7303_v = ~(v_w679_v | v_w1883_v);
	assign v_w2888_v = v_w552_v ^ v_w2887_v;
	assign v_w6198_v = ~(v_w1503_v | v_w6197_v);
	assign v_w2394_v = ~(v_w2357_v & v_s279_v);
	assign v_w363_v = ~(v_s502_v);
	assign v_w4841_v = ~(v_w1083_v | v_w2264_v);
	assign v_w1493_v = ~(v_w1051_v & v_s224_v);
	assign v_w5026_v = ~(v_w5018_v | v_w5025_v);
	assign v_w493_v = ~(v_w6646_v & v_w6653_v);
	assign v_w4455_v = ~(v_w1011_v & v_w2753_v);
	assign v_w1866_v = ~(v_w1094_v);
	assign v_w1472_v = ~(v_w1471_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s266_v<=0;
	end
	else
	begin
	v_s266_v<=v_w283_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s77_v<=0;
	end
	else
	begin
	v_s77_v<=v_w85_v;
	end
	end
	assign v_w6715_v = ~(v_w6714_v & v_w758_v);
	assign v_w5065_v = ~(v_w5064_v ^ v_w2459_v);
	assign v_w3210_v = ~(v_w3204_v & v_w3209_v);
	assign v_w1591_v = ~(v_w1590_v & v_w648_v);
	assign v_w3400_v = ~(v_s261_v & v_w3222_v);
	assign v_w531_v = ~(v_s520_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s64_v<=0;
	end
	else
	begin
	v_s64_v<=v_w72_v;
	end
	end
	assign v_w829_v = ~(v_w713_v | v_s268_v);
	assign v_w536_v = ~(v_w534_v | v_w535_v);
	assign v_w3512_v = ~(v_w3503_v | v_w3511_v);
	assign v_w4840_v = ~(v_w4838_v & v_w4839_v);
	assign v_w3001_v = ~(v_w2794_v | v_w3000_v);
	assign v_w808_v = ~(v_w672_v & v_w612_v);
	assign v_w1681_v = ~(v_w1445_v);
	assign v_w7056_v = ~(v_w7054_v & v_w7055_v);
	assign v_w5691_v = ~(v_w5689_v & v_w5690_v);
	assign v_w2539_v = ~(v_w2537_v | v_w2538_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s80_v<=0;
	end
	else
	begin
	v_s80_v<=v_w88_v;
	end
	end
	assign v_w3812_v = ~(v_w2847_v | v_w3735_v);
	assign v_w2329_v = ~(v_s172_v & v_s476_v);
	assign v_w6090_v = ~(v_w6088_v & v_w6089_v);
	assign v_w6547_v = ~(v_w6542_v | v_w888_v);
	assign v_w1045_v = ~(v_in17_v & v_w1229_v);
	assign v_w2024_v = ~(v_w986_v | v_w2023_v);
	assign v_w5840_v = ~(v_s287_v & v_w529_v);
	assign v_w299_v = ~(v_w4107_v & v_w4113_v);
	assign v_w3519_v = ~(v_w3518_v);
	assign v_w3649_v = ~(v_w3508_v | v_w3515_v);
	assign v_w4317_v = ~(v_w4316_v & v_w690_v);
	assign v_w2447_v = ~(v_w2284_v | v_w2242_v);
	assign v_w6322_v = ~(v_w6320_v & v_w6321_v);
	assign v_w8110_v = v_w6291_v & v_w6020_v;
	assign v_w411_v = ~(v_w7177_v & v_w7178_v);
	assign v_w6858_v = ~(v_w6857_v | v_w1684_v);
	assign v_w762_v = v_w2709_v & v_w2712_v;
	assign v_w2049_v = ~(v_w2046_v & v_w2048_v);
	assign v_w2933_v = ~(v_w2927_v | v_w2932_v);
	assign v_w7216_v = ~(v_w7117_v | v_w1517_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s237_v<=0;
	end
	else
	begin
	v_s237_v<=v_w250_v;
	end
	end
	assign v_w3996_v = ~(v_w871_v | v_w3731_v);
	assign v_w2208_v = ~(v_s155_v | v_s154_v);
	assign v_w3332_v = ~(v_w3109_v & v_w2429_v);
	assign v_w4228_v = ~(v_w4207_v & v_w4210_v);
	assign v_w5973_v = ~(v_w5971_v & v_w5972_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s68_v<=0;
	end
	else
	begin
	v_s68_v<=v_w76_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s341_v<=0;
	end
	else
	begin
	v_s341_v<=v_w374_v;
	end
	end
	assign v_w3348_v = ~(v_w760_v & v_w2639_v);
	assign v_w3428_v = ~(v_w3426_v | v_w3427_v);
	assign v_w7754_v = ~(v_w654_v & v_w7753_v);
	assign v_w2059_v = v_w1435_v | v_w2058_v;
	assign v_w144_v = v_s135_v & v_w5134_v;
	assign v_w3885_v = ~(v_w3883_v | v_w3884_v);
	assign v_w8_v = ~(v_s479_v);
	assign v_w756_v = ~(v_w755_v);
	assign v_w6177_v = ~(v_w6018_v | v_w1514_v);
	assign v_w7116_v = ~(v_w7114_v | v_w7115_v);
	assign v_w5514_v = ~(v_w4632_v & v_w5513_v);
	assign v_w2010_v = v_w1678_v & v_w2008_v;
	assign v_w2704_v = ~(v_w2701_v | v_w2703_v);
	assign v_w1318_v = ~(v_w1052_v & v_s31_v);
	assign v_w1555_v = ~(v_w713_v);
	assign v_w5924_v = ~(v_w5922_v & v_w5923_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s500_v<=0;
	end
	else
	begin
	v_s500_v<=v_w344_v;
	end
	end
	assign v_w402_v = ~(v_w3437_v & v_w3446_v);
	assign v_w5250_v = ~(v_w5248_v | v_w5249_v);
	assign v_w6037_v = ~(v_w6013_v & v_w6030_v);
	assign v_w6119_v = ~(v_w6029_v | v_w6118_v);
	assign v_w2100_v = ~(v_w2097_v & v_w1287_v);
	assign v_w2581_v = ~(v_s293_v ^ v_w2580_v);
	assign v_w5793_v = ~(v_s408_v & v_w529_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s363_v<=0;
	end
	else
	begin
	v_s363_v<=v_w406_v;
	end
	end
	assign v_w6427_v = ~(v_w6417_v & v_w6416_v);
	assign v_w1462_v = ~(v_w718_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s440_v<=0;
	end
	else
	begin
	v_s440_v<=v_w492_v;
	end
	end
	assign v_w7665_v = ~(v_w7664_v & v_w7097_v);
	assign v_w5154_v = ~(v_w5152_v | v_w5153_v);
	assign v_w4593_v = ~(v_w4592_v & v_w673_v);
	assign v_w1310_v = ~(v_w1065_v | v_w1309_v);
	assign v_w5743_v = ~(v_w5707_v & v_w1617_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s313_v<=0;
	end
	else
	begin
	v_s313_v<=v_w338_v;
	end
	end
	assign v_w3031_v = v_s380_v ^ v_w2651_v;
	assign v_w5479_v = ~(v_w683_v & v_w5478_v);
	assign v_w5728_v = ~(v_w1324_v | v_w2138_v);
	assign v_w2242_v = ~(v_w554_v & v_w2241_v);
	assign v_w805_v = ~(v_w803_v | v_w804_v);
	assign v_w3530_v = ~(v_w3525_v & v_w3529_v);
	assign v_w5916_v = v_w5915_v ^ v_w2070_v;
	assign v_w6039_v = ~(v_w6038_v & v_w533_v);
	assign v_w1641_v = ~(v_w1639_v & v_w1640_v);
	assign v_w7188_v = ~(v_w1467_v | v_w7117_v);
	assign v_w931_v = ~(v_w1814_v | v_w1882_v);
	assign v_w7489_v = ~(v_w7481_v & v_w7488_v);
	assign v_w5789_v = ~(v_w5787_v & v_w5788_v);
	assign v_w8034_v = ~(v_w7996_v | v_w8033_v);
	assign v_w5411_v = ~(v_w4863_v | v_w4855_v);
	assign v_w3656_v = ~(v_w3650_v | v_w3655_v);
	assign v_w3349_v = ~(v_w3347_v & v_w3348_v);
	assign v_w3183_v = ~(v_w625_v ^ v_w3182_v);
	assign v_w4143_v = ~(v_w4141_v & v_w4142_v);
	assign v_w4943_v = ~(v_w4940_v | v_w4942_v);
	assign v_w6755_v = ~(v_w6746_v & v_w6754_v);
	assign v_w3928_v = ~(v_w3783_v & v_w3780_v);
	assign v_w6997_v = ~(v_w884_v & v_w6996_v);
	assign v_w1402_v = ~(v_w847_v | v_w1401_v);
	assign v_w856_v = ~(v_w1111_v | v_w774_v);
	assign v_w7658_v = ~(v_w2105_v & v_w2129_v);
	assign v_w5843_v = ~(v_w2117_v & v_w1027_v);
	assign v_w4426_v = ~(v_w4397_v & v_w4425_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s109_v<=0;
	end
	else
	begin
	v_s109_v<=v_w117_v;
	end
	end
	assign v_w7822_v = ~(v_s417_v & v_w7742_v);
	assign v_w374_v = ~(v_w6853_v & v_w6869_v);
	assign v_w6933_v = ~(v_w6932_v & v_w1915_v);
	assign v_w242_v = ~(v_w5568_v & v_w5569_v);
	assign v_w4858_v = ~(v_w674_v & v_s364_v);
	assign v_w5431_v = ~(v_w5427_v | v_w5430_v);
	assign v_w713_v = v_s477_v | v_s265_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s34_v<=0;
	end
	else
	begin
	v_s34_v<=v_w38_v;
	end
	end
	assign v_w4639_v = ~(v_w4637_v | v_w4638_v);
	assign v_w5579_v = ~(v_w675_v & v_w5384_v);
	assign v_w5458_v = ~(v_w5123_v | v_w4741_v);
	assign v_w4583_v = ~(v_w3603_v & v_w4582_v);
	assign v_w1438_v = ~(v_w1436_v & v_w1437_v);
	assign v_w6854_v = ~(v_w1869_v ^ v_w1870_v);
	assign v_w1536_v = ~(v_w830_v & v_w944_v);
	assign v_w3630_v = ~(v_w3604_v & v_w873_v);
	assign v_w1780_v = ~(v_w1779_v | v_w8_v);
	assign v_w366_v = ~(v_w7189_v & v_w7190_v);
	assign v_w3911_v = ~(v_w3807_v & v_w3804_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s342_v<=0;
	end
	else
	begin
	v_s342_v<=v_w375_v;
	end
	end
	assign v_w4365_v = ~(v_w4363_v | v_w4364_v);
	assign v_w6975_v = ~(v_w6973_v & v_w6974_v);
	assign v_w5782_v = ~(v_w5774_v | v_w5781_v);
	assign v_w4940_v = ~(v_w4938_v & v_w4939_v);
	assign v_w264_v = ~(v_w5154_v & v_w5155_v);
	assign v_w5067_v = ~(v_w2448_v & v_w1131_v);
	assign v_w2910_v = ~(v_w2908_v & v_w2909_v);
	assign v_w2363_v = ~(v_w314_v ^ v_w2362_v);
	assign v_w7823_v = v_w8198_v ^ v_keyinput_94_v;
	assign v_w2702_v = ~(v_w432_v ^ v_w2656_v);
	assign v_w3566_v = ~(v_w3565_v);
	assign v_w5854_v = ~(v_w5852_v & v_w5853_v);
	assign v_w7419_v = ~(v_w7414_v & v_w7417_v);
	assign v_w5890_v = ~(v_w5888_v & v_w5889_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s403_v<=0;
	end
	else
	begin
	v_s403_v<=v_w452_v;
	end
	end
	assign v_w4852_v = ~(v_w4526_v | v_w4848_v);
	assign v_w3346_v = v_w3345_v ^ v_w3048_v;
	assign v_w2478_v = ~(v_w617_v);
	assign v_w3926_v = ~(v_w3791_v | v_w3925_v);
	assign v_w1956_v = ~(v_w1940_v | v_w1955_v);
	assign v_w2960_v = v_s162_v ^ v_w2959_v;
	assign v_w3833_v = ~(v_w2296_v & v_w3732_v);
	assign v_w7738_v = ~(v_w1096_v | v_w1782_v);
	assign v_w8095_v = ~(v_w2005_v | v_w2071_v);
	assign v_w4445_v = ~(v_w4444_v & v_w3485_v);
	assign v_w6291_v = ~(v_w6289_v ^ v_w6290_v);
	assign v_w3923_v = ~(v_w3921_v & v_w3922_v);
	assign v_w7883_v = ~(v_s114_v & v_w7876_v);
	assign v_w7609_v = ~(v_w1402_v | v_w7608_v);
	assign v_w601_v = ~(v_w2062_v | v_w2064_v);
	assign v_w4139_v = ~(v_w4138_v & v_w4130_v);
	assign v_w6101_v = ~(v_w6100_v & v_w6020_v);
	assign v_w3011_v = ~(v_w3009_v & v_w3010_v);
	assign v_w4816_v = ~(v_w4814_v | v_w4815_v);
	assign v_w4482_v = ~(v_w4480_v | v_w4481_v);
	assign v_w7346_v = ~(v_w1820_v | v_w680_v);
	assign v_w3874_v = v_w3868_v | v_w3865_v;
	assign v_w7932_v = ~(v_w527_v & v_w1135_v);
	assign v_w7490_v = v_w7487_v | v_w7484_v;
	assign v_w868_v = ~(v_w910_v & v_w911_v);
	assign v_w6679_v = v_w6678_v ^ v_w1744_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s96_v<=0;
	end
	else
	begin
	v_s96_v<=v_w104_v;
	end
	end
	assign v_w3237_v = ~(v_w3235_v | v_w3236_v);
	assign v_w3097_v = ~(v_w3088_v | v_w3096_v);
	assign v_w7205_v = ~(v_w7203_v | v_w7204_v);
	assign v_w7392_v = ~(v_w945_v | v_w680_v);
	assign v_w7430_v = ~(v_w7395_v & v_w7429_v);
	assign v_w2849_v = ~(v_s325_v & v_w565_v);
	assign v_w5813_v = ~(v_w892_v & v_w1095_v);
	assign v_w1560_v = ~(v_w615_v & v_s267_v);
	assign v_w1729_v = ~(v_w1119_v);
	assign v_w6912_v = v_w724_v | v_w1825_v;
	assign v_w6850_v = ~(v_w6848_v | v_w6849_v);
	assign v_w1777_v = ~(v_w685_v & v_w1776_v);
	assign v_w7484_v = ~(v_w7482_v | v_w7483_v);
	assign v_w7528_v = ~(v_w7524_v | v_w7527_v);
	assign v_w6002_v = ~(v_w1418_v | v_w2138_v);
	assign v_w2679_v = ~(v_w2677_v & v_w2678_v);
	assign v_w1066_v = ~(v_w1314_v & v_w1315_v);
	assign v_w3199_v = ~(v_w3195_v | v_w3198_v);
	assign v_w4390_v = ~(v_w4376_v & v_w4389_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s199_v<=0;
	end
	else
	begin
	v_s199_v<=v_w212_v;
	end
	end
	assign v_w837_v = ~(v_w1607_v | v_w808_v);
	assign v_w3276_v = ~(v_w3109_v & v_w2367_v);
	assign v_w5523_v = ~(v_w683_v & v_w5522_v);
	assign v_w5632_v = ~(v_s298_v & v_w695_v);
	assign v_w7295_v = ~(v_w680_v | v_w997_v);
	assign v_w2085_v = ~(v_w2082_v | v_w2084_v);
	assign v_w504_v = ~(v_w6581_v & v_w6582_v);
	assign v_w8200_v = v_w8199_v ^ v_keyinput_95_v;
	assign v_w796_v = ~(v_w794_v & v_w795_v);
	assign v_w399_v = ~(v_w3356_v & v_w3365_v);
	assign v_w2892_v = ~(v_w2889_v & v_w2891_v);
	assign v_w4407_v = ~(v_w2965_v | v_w4406_v);
	assign v_w5167_v = ~(v_w5146_v & v_w1299_v);
	assign v_w7933_v = ~(v_s208_v & v_w6015_v);
	assign v_w128_v = ~(v_w5582_v & v_w5583_v);
	assign v_w8098_v = ~(v_in27_v ^ v_w1262_v);
	assign v_w8047_v = ~(v_w7983_v | v_w8046_v);
	assign v_w6697_v = ~(v_w1798_v & v_w1323_v);
	assign v_w950_v = ~(v_w948_v | v_w949_v);
	assign v_w5456_v = ~(v_w5454_v | v_w5455_v);
	assign v_w19_v = ~(v_s480_v);
	assign v_w6901_v = ~(v_w6899_v & v_w6900_v);
	assign v_w3871_v = ~(v_w3859_v | v_w3856_v);
	assign v_w6338_v = ~(v_w6336_v | v_w6337_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s118_v<=0;
	end
	else
	begin
	v_s118_v<=v_w127_v;
	end
	end
	assign v_w84_v = ~(v_w7959_v & v_w7960_v);
	assign v_w1416_v = ~(v_w1414_v & v_w1415_v);
	assign v_w5644_v = ~(v_s193_v & v_w695_v);
	assign v_w2426_v = ~(v_w2422_v | v_w2425_v);
	assign v_w2193_v = v_s168_v ^ v_w2157_v;
	assign v_w1686_v = ~(v_w1680_v & v_w1685_v);
	assign v_w913_v = ~(v_w936_v | v_w1753_v);
	assign v_w7397_v = ~(v_w687_v | v_w578_v);
	assign v_w15_v = ~(v_w7971_v & v_w7972_v);
	assign v_w1934_v = ~(v_s70_v | v_s69_v);
	assign v_w629_v = v_w632_v | v_w633_v;
	assign v_w6414_v = ~(v_w1667_v & v_w6386_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s274_v<=0;
	end
	else
	begin
	v_s274_v<=v_w292_v;
	end
	end
	assign v_w7817_v = ~(v_w6660_v | v_w1919_v);
	assign v_w2408_v = ~(v_w8232_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s226_v<=0;
	end
	else
	begin
	v_s226_v<=v_w239_v;
	end
	end
	assign v_w5303_v = ~(v_w5109_v & v_w5302_v);
	assign v_w1791_v = ~(v_w1052_v & v_s9_v);
	assign v_w3296_v = ~(v_w3295_v & v_w3126_v);
	assign v_w1788_v = v_w1787_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s82_v<=0;
	end
	else
	begin
	v_s82_v<=v_w90_v;
	end
	end
	assign v_w6148_v = ~(v_w6018_v | v_w1528_v);
	assign v_w1963_v = ~(v_w1933_v | v_w1962_v);
	assign v_w3865_v = ~(v_w3863_v | v_w3864_v);
	assign v_w1871_v = ~(v_w1869_v & v_w1870_v);
	assign v_w925_v = ~(v_s327_v | v_s124_v);
	assign v_w2313_v = ~(v_w2312_v);
	assign v_w7636_v = ~(v_w6578_v);
	assign v_w1588_v = ~(v_w1548_v | v_w1587_v);
	assign v_w8239_v = v_w8238_v ^ v_keyinput_119_v;
	assign v_w6676_v = ~(v_w1067_v | v_w6579_v);
	assign v_w4223_v = ~(v_w3151_v | v_w4222_v);
	assign v_w184_v = ~(v_w5264_v & v_w5265_v);
	assign v_w421_v = ~(v_w4081_v & v_w4097_v);
	assign v_w3056_v = ~(v_s383_v ^ v_w2654_v);
	assign v_w1041_v = ~(v_w1062_v & v_s157_v);
	assign v_w8062_v = ~(v_w6113_v | v_w6117_v);
	assign v_w2903_v = ~(v_w2358_v & v_s331_v);
	assign v_w5989_v = ~(v_w662_v & v_w1309_v);
	assign v_w3262_v = ~(v_w872_v | v_w2620_v);
	assign v_w1661_v = ~(v_w1471_v | v_w1660_v);
	assign v_w3360_v = v_w3358_v ^ v_w3359_v;
	assign v_w3658_v = ~(v_w2383_v | v_w3657_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s458_v<=0;
	end
	else
	begin
	v_s458_v<=v_w511_v;
	end
	end
	assign v_w8196_v = ~(v_w783_v & v_w542_v);
	assign v_w3907_v = ~(v_w3899_v | v_w3906_v);
	assign v_w7620_v = ~(v_w7619_v & v_w1325_v);
	assign v_w5390_v = ~(v_w5388_v & v_w5389_v);
	assign v_w250_v = ~(v_w7923_v & v_w7924_v);
	assign v_w3260_v = ~(v_w3126_v & v_w3259_v);
	assign v_w6834_v = ~(v_w1428_v | v_w6571_v);
	assign v_w405_v = ~(v_w4887_v & v_w4897_v);
	assign v_w5998_v = ~(v_w5996_v | v_w5997_v);
	assign v_w3213_v = ~(v_w2639_v & v_w2803_v);
	assign v_w3386_v = ~(v_w3384_v ^ v_w3385_v);
	assign v_w7415_v = ~(v_w680_v | v_w1835_v);
	assign v_w6855_v = ~(v_w6854_v & v_w1915_v);
	assign v_w4024_v = ~(v_w4022_v & v_w4023_v);
	assign v_w5328_v = ~(v_w683_v & v_w5327_v);
	assign v_w5055_v = ~(v_w2343_v & v_w5054_v);
	assign v_w8225_v = ~(v_w5529_v | v_w5530_v);
	assign v_o17_v = v_w8004_v ^ v_w8013_v;
	assign v_w4945_v = ~(v_w4944_v & v_w2341_v);
	assign v_w4448_v = ~(v_w753_v & v_w2706_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s279_v<=0;
	end
	else
	begin
	v_s279_v<=v_w298_v;
	end
	end
	assign v_w960_v = ~(v_w778_v);
	assign v_w5015_v = ~(v_w5013_v | v_w5014_v);
	assign v_w3221_v = v_w2626_v & v_w2633_v;
	assign v_w7105_v = ~(v_w655_v & v_w7104_v);
	assign v_w5051_v = ~(v_w5049_v & v_w5050_v);
	assign v_w6115_v = ~(v_w657_v & v_s273_v);
	assign v_w2122_v = ~(v_w2120_v | v_w2121_v);
	assign v_w2522_v = ~(v_w2520_v & v_w2521_v);
	assign v_w24_v = ~(v_w7967_v & v_w7968_v);
	assign v_w8198_v = ~(v_w962_v | v_w1782_v);
	assign v_w5446_v = ~(v_w8157_v);
	assign v_w4770_v = ~(v_w4526_v | v_w4766_v);
	assign v_w342_v = ~(v_w4220_v & v_w4221_v);
	assign v_w5694_v = ~(v_w728_v ^ v_w2031_v);
	assign v_w7094_v = ~(v_w7092_v & v_w7093_v);
	assign v_w1159_v = ~(v_s342_v | v_w1158_v);
	assign v_w2828_v = ~(v_w2827_v | v_w617_v);
	assign v_w8011_v = v_s377_v ^ v_s456_v;
	assign v_w8145_v = v_w8144_v ^ v_keyinput_55_v;
	assign v_w1226_v = ~(v_w1224_v & v_w1225_v);
	assign v_w3164_v = ~(v_w2607_v & v_w1131_v);
	assign v_w7762_v = ~(v_w1020_v | v_w1782_v);
	assign v_w3388_v = ~(v_w2901_v & v_w2639_v);
	assign v_w4592_v = ~(v_w4532_v & v_w4591_v);
	assign v_w5439_v = ~(v_w5437_v & v_w5438_v);
	assign v_w393_v = ~(v_w6801_v & v_w6817_v);
	assign v_w6789_v = v_w758_v & v_w6787_v;
	assign v_w571_v = ~(v_w1467_v | v_w2294_v);
	assign v_w3767_v = v_w3763_v | v_w3766_v;
	assign v_w1610_v = ~(v_s319_v ^ v_w1609_v);
	assign v_w5198_v = ~(v_w5196_v | v_w5197_v);
	assign v_w4_v = ~(v_w7977_v & v_w7978_v);
	assign v_w3052_v = ~(v_w2478_v & v_w851_v);
	assign v_w7644_v = ~(v_w7557_v & v_w7643_v);
	assign v_w3477_v = v_w855_v ^ v_w3460_v;
	assign v_w4391_v = ~(v_w4390_v ^ v_s394_v);
	assign v_w5723_v = ~(v_w1337_v ^ v_w2083_v);
	assign v_w6500_v = ~(v_s355_v ^ v_w6499_v);
	assign v_w7013_v = ~(v_s288_v & v_w656_v);
	assign v_w1435_v = ~(v_w1433_v & v_w1434_v);
	assign v_w161_v = v_s152_v & v_w5134_v;
	assign v_w5308_v = ~(v_w5124_v & v_w5085_v);
	assign v_w4648_v = ~(v_w4647_v & v_w878_v);
	assign v_w5715_v = ~(v_w5713_v & v_w5714_v);
	assign v_w7690_v = ~(v_w7042_v & v_w7689_v);
	assign v_w2881_v = ~(v_s347_v | v_w2880_v);
	assign v_w7763_v = ~(v_w6827_v | v_w7762_v);
	assign v_w1863_v = ~(v_w1822_v & v_w1862_v);
	assign v_w7373_v = ~(v_w687_v | v_w989_v);
	assign v_w7442_v = ~(v_w7440_v | v_w7441_v);
	assign v_w1954_v = ~(v_w1950_v | v_w1953_v);
	assign v_w125_v = ~(v_w5588_v & v_w5589_v);
	assign v_w5132_v = ~(v_w674_v | v_w5131_v);
	assign v_w3243_v = ~(v_w2940_v | v_w2943_v);
	assign v_w870_v = ~(v_w667_v | v_w730_v);
	assign v_w2845_v = ~(v_w699_v & v_s201_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s423_v<=0;
	end
	else
	begin
	v_s423_v<=v_w474_v;
	end
	end
	assign v_w7737_v = ~(v_w6894_v | v_w1919_v);
	assign v_w1923_v = ~(v_w1921_v & v_w1922_v);
	assign v_w203_v = ~(v_w5534_v & v_w5541_v);
	assign v_w3734_v = ~(v_w1068_v | v_w3731_v);
	assign v_w65_v = v_s57_v & v_w7107_v;
	assign v_w7000_v = ~(v_w6996_v & v_w758_v);
	assign v_w1386_v = v_w746_v ^ v_w747_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s491_v<=0;
	end
	else
	begin
	v_s491_v<=v_w265_v;
	end
	end
	assign v_w5879_v = ~(v_w662_v & v_w578_v);
	assign v_w3916_v = ~(v_w3915_v & v_w881_v);
	assign v_w2326_v = v_w2324_v & v_w2325_v;
	assign v_w1302_v = v_s438_v ^ v_w1168_v;
	assign v_w5920_v = ~(v_w1718_v | v_w2135_v);
	assign v_w3022_v = v_w552_v ^ v_w3021_v;
	assign v_w6166_v = ~(v_w1528_v | v_w6144_v);
	assign v_w6003_v = ~(v_w6001_v | v_w6002_v);
	assign v_w2737_v = ~(v_w2355_v & v_s94_v);
	assign v_w2798_v = v_w531_v & v_s217_v;
	assign v_w3518_v = ~(v_w2803_v | v_w2619_v);
	assign v_w2846_v = ~(v_w2844_v & v_w2845_v);
	assign v_w2669_v = ~(v_w2666_v | v_w2668_v);
	assign v_w7224_v = ~(v_w7117_v | v_w1542_v);
	assign v_w1_v = ~(v_s478_v);
	assign v_w5207_v = ~(v_s115_v & v_w5141_v);
	assign v_w2552_v = ~(v_s291_v | v_w2551_v);
	assign v_w6380_v = ~(v_w6351_v | v_w6355_v);
	assign v_w2035_v = ~(v_w723_v ^ v_w839_v);
	assign v_w993_v = ~(v_w992_v);
	assign v_w3207_v = ~(v_w3109_v & v_w2833_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s186_v<=0;
	end
	else
	begin
	v_s186_v<=v_w199_v;
	end
	end
	assign v_w5013_v = v_s296_v & v_w674_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s38_v<=0;
	end
	else
	begin
	v_s38_v<=v_w45_v;
	end
	end
	assign v_w6457_v = ~(v_w1407_v);
	assign v_w5302_v = ~(v_w5098_v | v_w5301_v);
	assign v_w1442_v = ~(v_w1439_v & v_w1441_v);
	assign v_w6255_v = ~(v_w1474_v ^ v_w6254_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s240_v<=0;
	end
	else
	begin
	v_s240_v<=v_w253_v;
	end
	end
	assign v_w5462_v = ~(v_s183_v & v_w5386_v);
	assign v_w1138_v = ~(v_w2242_v & v_w2602_v);
	assign v_w1764_v = ~(v_s11_v & v_w1103_v);
	assign v_w850_v = ~(v_w848_v | v_w849_v);
	assign v_w5060_v = ~(v_s277_v | v_w2261_v);
	assign v_w2850_v = ~(v_w2777_v | v_w531_v);
	assign v_w3657_v = ~(v_w3648_v & v_w3656_v);
	assign v_w3948_v = ~(v_w3735_v & v_w3558_v);
	assign v_w4171_v = ~(v_w2604_v & v_w4170_v);
	assign v_w398_v = ~(v_w7854_v & v_w7855_v);
	assign v_w2266_v = ~(v_w1136_v);
	assign v_w2885_v = ~(v_w2884_v & v_w569_v);
	assign v_w1543_v = ~(v_w1542_v | v_w808_v);
	assign v_w4716_v = ~(v_w2265_v & v_w820_v);
	assign v_w3965_v = ~(v_w3957_v | v_w3964_v);
	assign v_w2430_v = ~(v_w2331_v | v_w2429_v);
	assign v_w4161_v = ~(v_w2290_v & v_s231_v);
	assign v_w351_v = ~(v_w7935_v & v_w7936_v);
	assign v_w5007_v = v_w3650_v ^ v_w4465_v;
	assign v_w6974_v = ~(v_w1140_v & v_w1484_v);
	assign v_w8192_v = v_w8191_v ^ v_keyinput_90_v;
	assign v_w7138_v = ~(v_w7136_v | v_w7137_v);
	assign v_w2192_v = ~(v_w2164_v & v_w2191_v);
	assign v_w5846_v = ~(v_w5842_v | v_w5845_v);
	assign v_w7518_v = ~(v_w7516_v & v_w7517_v);
	assign v_w2_v = ~(v_w5685_v);
	assign v_w182_v = ~(v_w5186_v & v_w5187_v);
	assign v_w4996_v = ~(v_w4863_v | v_w4995_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s257_v<=0;
	end
	else
	begin
	v_s257_v<=v_w272_v;
	end
	end
	assign v_w5295_v = ~(v_w2258_v & v_w2419_v);
	assign v_w5050_v = ~(v_w2384_v & v_w2347_v);
	assign v_w2564_v = ~(v_w2561_v | v_w2563_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s356_v<=0;
	end
	else
	begin
	v_s356_v<=v_w394_v;
	end
	end
	assign v_w5816_v = ~(v_w1459_v & v_w5707_v);
	assign v_w4175_v = ~(v_w4160_v & v_w4163_v);
	assign v_w5935_v = ~(v_w5934_v & v_w5703_v);
	assign v_w1917_v = ~(v_w1802_v & v_w1916_v);
	assign v_w2724_v = ~(v_w2714_v & v_w2723_v);
	assign v_w4375_v = ~(v_w4371_v | v_w4374_v);
	assign v_w2854_v = ~(v_w2849_v & v_w2853_v);
	assign v_w36_v = ~(v_w7963_v & v_w7964_v);
	assign v_w977_v = ~(v_in25_v ^ v_w1255_v);
	assign v_w7365_v = ~(v_w7360_v & v_w7363_v);
	assign v_w4282_v = ~(v_w4281_v & v_w690_v);
	assign v_w8076_v = v_w8075_v ^ v_keyinput_11_v;
	assign v_w3770_v = ~(v_w3768_v & v_w3769_v);
	assign v_w8170_v = v_w8169_v ^ v_keyinput_74_v;
	assign v_w5981_v = ~(v_w892_v & v_w789_v);
	assign v_w6658_v = ~(v_w6656_v | v_w6657_v);
	assign v_w5987_v = ~(v_w5985_v | v_w5986_v);
	assign v_w3606_v = ~(v_w3605_v & v_w3595_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s520_v<=0;
	end
	else
	begin
	v_s520_v<=v_w530_v;
	end
	end
	assign v_w5868_v = ~(v_w1311_v | v_w2138_v);
	assign v_w2379_v = ~(v_w2378_v);
	assign v_w1039_v = ~(v_w8236_v);
	assign v_w5874_v = ~(v_w1316_v | v_w2135_v);
	assign v_w6062_v = ~(v_w6060_v & v_w6061_v);
	assign v_w3196_v = ~(v_w699_v & v_s190_v);
	assign v_w274_v = ~(v_s492_v);
	assign v_w1168_v = v_w1167_v | v_s436_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s484_v<=0;
	end
	else
	begin
	v_s484_v<=v_w41_v;
	end
	end
	assign v_w6396_v = ~(v_w1667_v & v_w6372_v);
	assign v_w6675_v = ~(v_w6673_v & v_w6674_v);
	assign v_w5228_v = ~(v_w693_v | v_w2822_v);
	assign v_w4611_v = ~(v_w4606_v & v_w4610_v);
	assign v_w4876_v = ~(v_w4874_v & v_w4875_v);
	assign v_w2520_v = ~(v_w2511_v & v_w2519_v);
	assign v_w6717_v = ~(v_w6710_v | v_w6716_v);
	assign v_w6835_v = v_w656_v & v_s354_v;
	assign v_w8166_v = v_w3853_v | v_w3876_v;
	assign v_w1716_v = ~(v_w1715_v & v_w809_v);
	assign v_w5735_v = ~(v_w1856_v | v_w5734_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s107_v<=0;
	end
	else
	begin
	v_s107_v<=v_w115_v;
	end
	end
	assign v_w6128_v = v_s286_v ^ v_w1528_v;
	assign v_w422_v = ~(v_w4125_v & v_w4134_v);
	assign v_w7947_v = ~(v_s90_v & v_w2143_v);
	assign v_w7398_v = ~(v_w7396_v | v_w7397_v);
	assign v_w645_v = ~(v_w981_v);
	assign v_w5797_v = ~(v_w5795_v | v_w5796_v);
	assign v_w6773_v = ~(v_w6764_v | v_w6772_v);
	assign v_w5340_v = ~(v_w5016_v & v_w5339_v);
	assign v_w2940_v = v_w2934_v & v_w2939_v;
	assign v_w2576_v = ~(v_w558_v & v_w2575_v);
	assign v_w650_v = ~(v_w1975_v & v_w1991_v);
	assign v_w7520_v = ~(v_w7518_v & v_w7519_v);
	assign v_w7811_v = v_w8209_v ^ v_keyinput_101_v;
	assign v_w8119_v = v_w575_v ^ v_keyinput_40_v;
	assign v_w5116_v = ~(v_s262_v & v_w674_v);
	assign v_w2636_v = ~(v_w8131_v);
	assign v_w2816_v = ~(v_w2815_v & v_w697_v);
	assign v_w9_v = ~(v_w7975_v & v_w7976_v);
	assign v_w3548_v = ~(v_w3544_v & v_w3547_v);
	assign v_w560_v = ~(v_s2_v | v_w559_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s307_v<=0;
	end
	else
	begin
	v_s307_v<=v_w330_v;
	end
	end
	assign v_w5094_v = ~(v_w5091_v | v_w5093_v);
	assign v_w3533_v = ~(v_w3531_v | v_w3532_v);
	assign v_w5799_v = v_w2072_v ^ v_w5798_v;
	assign v_w1537_v = ~(v_s242_v & v_w561_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s187_v<=0;
	end
	else
	begin
	v_s187_v<=v_w200_v;
	end
	end
	assign v_w2551_v = v_w531_v | v_w2550_v;
	assign v_w5354_v = ~(v_s211_v & v_w5293_v);
	assign v_w3364_v = ~(v_w3121_v | v_w825_v);
	assign v_w2219_v = ~(v_w2215_v | v_w2218_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s483_v<=0;
	end
	else
	begin
	v_s483_v<=v_w39_v;
	end
	end
	assign v_w7557_v = ~(v_w7556_v & v_w1775_v);
	assign v_w7962_v = ~(v_w527_v & v_w1337_v);
	assign v_w7803_v = ~(v_s75_v & v_w7742_v);
	assign v_w1193_v = ~(v_s18_v & v_w1192_v);
	assign v_w6662_v = ~(v_w6661_v & v_w884_v);
	assign v_w8007_v = v_w280_v & v_w8006_v;
	assign v_w482_v = ~(v_w5670_v & v_w5671_v);
	assign v_w2984_v = v_w384_v ^ v_w2983_v;
	assign v_w1627_v = ~(v_w1374_v | v_w1626_v);
	assign v_w4814_v = ~(v_w4812_v & v_w4813_v);
	assign v_w2044_v = ~(v_w2032_v & v_w1135_v);
	assign v_w5827_v = ~(v_w5825_v | v_w5826_v);
	assign v_w2825_v = ~(v_w2821_v & v_w2824_v);
	assign v_w4968_v = ~(v_w4967_v & v_w878_v);
	assign v_w6579_v = ~(v_w2126_v & v_w1141_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s366_v<=0;
	end
	else
	begin
	v_s366_v<=v_w409_v;
	end
	end
	assign v_w4081_v = ~(v_w4072_v | v_w4080_v);
	assign v_w6412_v = ~(v_w6408_v ^ v_w6411_v);
	assign v_w2967_v = ~(v_w2956_v);
	assign v_w7204_v = ~(v_w1476_v | v_w7117_v);
	assign v_w3553_v = ~(v_w2791_v & v_w967_v);
	assign v_w2560_v = v_w2548_v & v_w2559_v;
	assign v_w1779_v = ~(v_s96_v | v_w1773_v);
	assign v_w6767_v = ~(v_w1814_v | v_w932_v);
	assign v_w2457_v = ~(v_w2456_v);
	assign v_w4148_v = ~(v_w4146_v & v_w4147_v);
	assign v_w6512_v = ~(v_w6490_v & v_w6493_v);
	assign v_w272_v = ~(v_w5294_v & v_w5297_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s448_v<=0;
	end
	else
	begin
	v_s448_v<=v_w501_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s192_v<=0;
	end
	else
	begin
	v_s192_v<=v_w205_v;
	end
	end
	assign v_w4470_v = ~(v_w8239_v);
	assign v_w7560_v = ~(v_w7558_v & v_w7559_v);
	assign v_w1071_v = ~(v_w1406_v & v_w1408_v);
	assign v_w2046_v = ~(v_w2038_v & v_w905_v);
	assign v_w3643_v = ~(v_w3642_v);
	assign v_w2648_v = ~(v_w2647_v & v_s361_v);
	assign v_w714_v = ~(v_w588_v & v_w324_v);
	assign v_w4451_v = ~(v_w760_v & v_w2738_v);
	assign v_w3796_v = ~(v_w3795_v & v_w2956_v);
	assign v_w1099_v = ~(v_w1097_v | v_w1098_v);
	assign v_w6849_v = ~(v_w1091_v | v_w6579_v);
	assign v_w6628_v = ~(v_w6624_v & v_w6627_v);
	assign v_w4958_v = ~(v_w2827_v | v_w2264_v);
	assign v_w709_v = ~(v_w2149_v | v_w2152_v);
	assign v_w2435_v = ~(v_w2434_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s209_v<=0;
	end
	else
	begin
	v_s209_v<=v_w222_v;
	end
	end
	assign v_w4607_v = ~(v_w4581_v & v_w873_v);
	assign v_w8030_v = ~(v_w7998_v | v_w8029_v);
	assign v_w238_v = ~(v_w7704_v & v_w7705_v);
	assign v_w66_v = v_s58_v & v_w7107_v;
	assign v_w5386_v = ~(v_w683_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s362_v<=0;
	end
	else
	begin
	v_s362_v<=v_w405_v;
	end
	end
	assign v_w2917_v = ~(v_w2916_v | v_w538_v);
	assign v_w7526_v = ~(v_w680_v & v_w961_v);
	assign v_w6159_v = ~(v_w6131_v & v_w6134_v);
	assign v_w792_v = ~(v_s173_v | v_w2154_v);
	assign v_w4708_v = ~(v_w4701_v & v_w4707_v);
	assign v_w5967_v = ~(v_w1373_v | v_w2138_v);
	assign v_w3252_v = ~(v_w3250_v | v_w3251_v);
	assign v_w7201_v = ~(v_w7199_v | v_w7200_v);
	assign v_w4707_v = ~(v_w4704_v | v_w4706_v);
	assign v_w4624_v = ~(v_w4621_v | v_w4623_v);
	assign v_w7141_v = v_w7113_v & v_s423_v;
	assign v_w1719_v = ~(v_w1718_v | v_w1180_v);
	assign v_w963_v = ~(v_w1120_v & v_w1121_v);
	assign v_w6319_v = ~(v_w6318_v & v_w659_v);
	assign v_w7115_v = ~(v_w528_v | v_w667_v);
	assign v_w3912_v = ~(v_w3910_v & v_w3911_v);
	assign v_w1259_v = v_in26_v ^ v_w1258_v;
	assign v_w2880_v = ~(v_w2879_v | v_w531_v);
	assign v_w4952_v = ~(v_w4950_v & v_w4951_v);
	assign v_w451_v = ~(v_w6780_v & v_w6781_v);
	assign v_w7694_v = ~(v_w7693_v | v_w7016_v);
	assign v_w2777_v = ~(v_s312_v | v_w2776_v);
	assign v_w6644_v = ~(v_w6592_v & v_w961_v);
	assign v_w2405_v = v_w2357_v & v_s266_v;
	assign v_w82_v = v_s74_v & v_w7107_v;
	assign v_w3311_v = ~(v_w3309_v | v_w3310_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s230_v<=0;
	end
	else
	begin
	v_s230_v<=v_w243_v;
	end
	end
	assign v_w1087_v = ~(v_w1443_v | v_w2294_v);
	assign v_w2042_v = v_w1606_v & v_w2035_v;
	assign v_w4191_v = ~(v_w4190_v ^ v_s212_v);
	assign v_w2120_v = ~(v_w2118_v & v_w2119_v);
	assign v_w741_v = ~(v_w8099_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s249_v<=0;
	end
	else
	begin
	v_s249_v<=v_w262_v;
	end
	end
	assign v_w4166_v = ~(v_w4159_v & v_w4165_v);
	assign v_w1051_v = ~(v_w668_v | v_w730_v);
	assign v_w6497_v = ~(v_w6458_v & v_w6456_v);
	assign v_w1642_v = ~(v_w1637_v | v_w1641_v);
	assign v_w3182_v = ~(v_w3045_v & v_w3047_v);
	assign v_w2805_v = ~(v_w558_v & v_w2618_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s44_v<=0;
	end
	else
	begin
	v_s44_v<=v_w52_v;
	end
	end
	assign v_w6805_v = ~(v_w6595_v & v_w6804_v);
	assign v_w6949_v = ~(v_w6595_v & v_w6948_v);
	assign v_w6422_v = ~(v_w6420_v & v_w6421_v);
	assign v_w6311_v = ~(v_w6309_v | v_w6310_v);
	assign v_w3752_v = ~(v_w881_v | v_w3597_v);
	assign v_w6922_v = ~(v_w6916_v ^ v_w726_v);
	assign v_w6963_v = ~(v_w1852_v ^ v_w6962_v);
	assign v_w3279_v = ~(v_w3278_v & v_w3126_v);
	assign v_w3046_v = ~(v_w625_v & v_w3045_v);
	assign v_w4861_v = ~(v_w1088_v | v_w2264_v);
	assign v_w4878_v = ~(v_w4866_v & v_w4877_v);
	assign v_w775_v = ~(v_s248_v & v_w1192_v);
	assign v_w2255_v = ~(v_w2253_v | v_w2254_v);
	assign v_w7167_v = ~(v_w1391_v | v_w529_v);
	assign v_w6206_v = v_w8172_v ^ v_keyinput_76_v;
	assign v_w1784_v = ~(v_w679_v | v_w1783_v);
	assign v_w6287_v = ~(v_w1610_v & v_w6262_v);
	assign v_w898_v = ~(v_w568_v);
	assign v_w1857_v = ~(v_w1856_v & v_w839_v);
	assign v_w7569_v = ~(v_w1661_v & v_w7568_v);
	assign v_w8169_v = ~(v_w5172_v | v_w5173_v);
	assign v_w5442_v = ~(v_w4783_v & v_w5441_v);
	assign v_w5484_v = ~(v_w4685_v | v_w5123_v);
	assign v_w4775_v = ~(v_w4772_v | v_w4774_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s112_v<=0;
	end
	else
	begin
	v_s112_v<=v_w121_v;
	end
	end
	assign v_w5187_v = ~(v_w8092_v);
	assign v_w3615_v = ~(v_w3489_v & v_w3614_v);
	assign v_w1260_v = ~(v_s227_v & v_w1103_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s89_v<=0;
	end
	else
	begin
	v_s89_v<=v_w97_v;
	end
	end
	assign v_w4817_v = ~(v_w415_v | v_w673_v);
	assign v_w4075_v = ~(v_w4067_v & v_w4044_v);
	assign v_w437_v = ~(v_s515_v);
	assign v_w6404_v = ~(v_w657_v & v_s341_v);
	assign v_w6452_v = ~(v_w6447_v & v_w6451_v);
	assign v_w8183_v = v_w1751_v & v_w1752_v;
	assign v_w7075_v = ~(v_w1788_v & v_w1834_v);
	assign v_w2820_v = ~(v_w2819_v | v_w538_v);
	assign v_w3406_v = ~(v_w3404_v & v_w3405_v);
	assign v_w7928_v = ~(v_w527_v & v_w788_v);
	assign v_w6302_v = ~(v_w1610_v & v_w6277_v);
	assign v_w5912_v = ~(v_w5910_v & v_w5911_v);
	assign v_w5416_v = ~(v_w5413_v & v_w5415_v);
	assign v_w5492_v = ~(v_w5037_v & v_w4673_v);
	assign v_w642_v = v_w1828_v ^ v_w2011_v;
	assign v_w3978_v = ~(v_w3974_v | v_w3977_v);
	assign v_w707_v = v_w705_v & v_w706_v;
	assign v_w4898_v = v_s350_v & v_w674_v;
	assign v_w5659_v = ~(v_w420_v & v_w3338_v);
	assign v_w1908_v = ~(v_w1805_v | v_w1907_v);
	assign v_w555_v = ~(v_w2233_v);
	assign v_w8128_v = v_w8127_v ^ v_keyinput_45_v;
	assign v_w4118_v = ~(v_w2312_v & v_s279_v);
	assign v_w6740_v = ~(v_w6738_v | v_w6739_v);
	assign v_w1257_v = ~(v_w612_v & v_s222_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s404_v<=0;
	end
	else
	begin
	v_s404_v<=v_w453_v;
	end
	end
	assign v_w5457_v = ~(v_w4749_v);
	assign v_w6631_v = ~(v_w758_v & v_w6619_v);
	assign v_w5896_v = ~(v_w2033_v & v_w5776_v);
	assign v_w8006_v = ~(v_s259_v & v_s454_v);
	assign v_w5382_v = ~(v_w4926_v | v_w5123_v);
	assign v_w6189_v = ~(v_s234_v & v_w6161_v);
	assign v_w3488_v = ~(v_w3485_v | v_w1069_v);
	assign v_w8059_v = ~(v_w7991_v | v_w7992_v);
	assign v_w8125_v = ~(v_w4318_v & v_w4304_v);
	assign v_w4549_v = ~(v_w3535_v & v_w4548_v);
	assign v_w7577_v = ~(v_w6767_v | v_w799_v);
	assign v_w6957_v = ~(v_w758_v & v_w6948_v);
	assign v_w3156_v = ~(v_w3150_v & v_w3155_v);
	assign v_w4743_v = ~(v_w2369_v & v_w2722_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s262_v<=0;
	end
	else
	begin
	v_s262_v<=v_w278_v;
	end
	end
	assign v_w1601_v = ~(v_w1599_v & v_w1600_v);
	assign v_w5732_v = ~(v_w5730_v | v_w5731_v);
	assign v_w6645_v = ~(v_w6643_v & v_w6644_v);
	assign v_w5436_v = ~(v_w864_v | v_w2602_v);
	assign v_w7073_v = ~(v_w7069_v & v_w758_v);
	assign v_w7313_v = ~(v_w7311_v | v_w7312_v);
	assign v_w7632_v = ~(v_w6569_v | v_w1796_v);
	assign v_w2937_v = ~(v_w2926_v);
	assign v_w7570_v = ~(v_w7567_v | v_w7569_v);
	assign v_w5613_v = ~(v_w5555_v & v_w5532_v);
	assign v_w5451_v = ~(v_w683_v & v_w5450_v);
	assign v_w2148_v = ~(v_w926_v);
	assign v_w5818_v = ~(v_w662_v & v_w1323_v);
	assign v_w83_v = ~(v_w7802_v & v_w7803_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s67_v<=0;
	end
	else
	begin
	v_s67_v<=v_w75_v;
	end
	end
	assign v_w1914_v = ~(v_w685_v & v_w1772_v);
	assign v_w5502_v = ~(v_w5037_v & v_w4645_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s468_v<=0;
	end
	else
	begin
	v_s468_v<=v_w521_v;
	end
	end
	assign v_w4802_v = ~(v_w4798_v | v_w4801_v);
	assign v_w5294_v = ~(v_s257_v & v_w5293_v);
	assign v_w6173_v = v_w1514_v | v_w6171_v;
	assign v_w6323_v = ~(v_s197_v & v_w888_v);
	assign v_w4752_v = ~(v_w674_v | v_w4751_v);
	assign v_w611_v = ~(v_w609_v | v_w610_v);
	assign v_w4867_v = v_w958_v ^ v_w4485_v;
	assign v_w3329_v = ~(v_w1099_v ^ v_w2836_v);
	assign v_w5469_v = ~(v_w4729_v | v_w5468_v);
	assign v_w1242_v = ~(v_w1240_v & v_w1241_v);
	assign v_w3459_v = ~(v_w3457_v & v_w3458_v);
	assign v_w523_v = ~(v_w6460_v & v_w6480_v);
	assign v_w2163_v = ~(v_s165_v ^ v_w2159_v);
	assign v_w1264_v = ~(v_w612_v & v_s232_v);
	assign v_w5362_v = ~(v_s209_v & v_w5293_v);
	assign v_w6453_v = ~(v_w6441_v | v_w6452_v);
	assign v_w1685_v = ~(v_w1683_v | v_w1684_v);
	assign v_w3869_v = ~(v_w3865_v & v_w3868_v);
	assign v_w3205_v = ~(v_s1_v | v_w337_v);
	assign v_w3317_v = ~(v_w2384_v & v_w2634_v);
	assign v_w1239_v = v_in20_v ^ v_w1238_v;
	assign v_w4221_v = ~(v_w2823_v & v_w887_v);
	assign v_w6941_v = ~(v_w6939_v & v_w6940_v);
	assign v_w2336_v = ~(v_w2331_v & v_w2335_v);
	assign v_w3904_v = ~(v_w2901_v & v_w881_v);
	assign v_w2403_v = ~(v_s253_v & v_w593_v);
	assign v_w2134_v = ~(v_w528_v | v_w2133_v);
	assign v_w2206_v = ~(v_w2204_v & v_w2205_v);
	assign v_w1890_v = ~(v_w1736_v & v_w1889_v);
	assign v_w6241_v = v_s215_v ^ v_w1474_v;
	assign v_w6562_v = ~(v_w6557_v & v_w6561_v);
	assign v_w7907_v = ~(v_s447_v & v_w1993_v);
	assign v_w5672_v = ~(v_s34_v & v_w695_v);
	assign v_w5160_v = v_w2191_v & v_s1_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s111_v<=0;
	end
	else
	begin
	v_s111_v<=v_w119_v;
	end
	end
	assign v_w6260_v = ~(v_s308_v & v_w1474_v);
	assign v_w7832_v = ~(v_w1783_v & v_w1003_v);
	assign v_w6235_v = ~(v_w1490_v & v_w6217_v);
	assign v_w2456_v = ~(v_w553_v | v_w2455_v);
	assign v_w4096_v = ~(v_w4094_v | v_w4095_v);
	assign v_w1299_v = ~(v_w842_v ^ v_w1058_v);
	assign v_w1707_v = ~(v_w1699_v & v_w1074_v);
	assign v_w2555_v = ~(v_w2554_v | v_w568_v);
	assign v_w3762_v = ~(v_w851_v & v_w881_v);
	assign v_w1483_v = ~(v_w874_v & v_s308_v);
	assign v_w6099_v = v_w1539_v ^ v_w6098_v;
	assign v_w1747_v = ~(v_w1312_v | v_w1746_v);
	assign v_w7348_v = v_w7344_v | v_w7347_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s297_v<=0;
	end
	else
	begin
	v_s297_v<=v_w319_v;
	end
	end
	assign v_w7124_v = ~(v_w890_v | v_w529_v);
	assign v_w1802_v = ~(v_w1790_v | v_w1801_v);
	assign v_w4744_v = ~(v_w3633_v ^ v_w4566_v);
	assign v_w4216_v = ~(v_w4214_v | v_w4215_v);
	assign v_w4837_v = ~(v_w4836_v & v_w673_v);
	assign v_w3313_v = ~(v_w3109_v & v_w2379_v);
	assign v_w773_v = ~(v_in5_v ^ v_w1276_v);
	assign v_w3192_v = ~(v_w3113_v | v_w437_v);
	assign v_w5082_v = ~(v_w5081_v & v_w878_v);
	assign v_w1214_v = v_in12_v ^ v_w1213_v;
	assign v_w6904_v = ~(v_w656_v | v_w6903_v);
	assign v_w2340_v = v_w2339_v ^ v_w2296_v;
	assign v_w4516_v = ~(v_w2690_v | v_w755_v);
	assign v_w3569_v = ~(v_w761_v & v_w2738_v);
	assign v_w3214_v = ~(v_w2505_v ^ v_w2508_v);
	assign v_w4929_v = ~(v_w4922_v & v_w4928_v);
	assign v_w3830_v = ~(v_w3735_v & v_w2379_v);
	assign v_w3098_v = ~(v_w3087_v);
	assign v_w1720_v = ~(v_w666_v & v_s91_v);
	assign v_w6434_v = ~(v_s114_v & v_w888_v);
	assign v_w7071_v = ~(v_w603_v ^ v_w1840_v);
	assign v_w5415_v = ~(v_w5414_v | v_w4851_v);
	assign v_w6813_v = ~(v_w1798_v & v_w895_v);
	assign v_w5423_v = ~(v_w5419_v | v_w5422_v);
	assign v_w3803_v = ~(v_w881_v | v_w2935_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s424_v<=0;
	end
	else
	begin
	v_s424_v<=v_w475_v;
	end
	end
	assign v_w7369_v = ~(v_w680_v | v_w766_v);
	assign v_w3899_v = ~(v_w3897_v & v_w3898_v);
	assign v_w3891_v = ~(v_w3829_v & v_w3890_v);
	assign v_w4638_v = ~(v_w2261_v | v_w2686_v);
	assign v_w5805_v = ~(v_w1642_v | v_w5734_v);
	assign v_w1653_v = ~(v_w1651_v | v_w1652_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s304_v<=0;
	end
	else
	begin
	v_s304_v<=v_w327_v;
	end
	end
	assign v_w6141_v = ~(v_w6139_v | v_w6140_v);
	assign v_w7612_v = ~(v_w1712_v | v_w7611_v);
	assign v_w1741_v = ~(v_w1338_v & v_w1740_v);
	assign v_w6237_v = ~(v_w6235_v & v_w6236_v);
	assign v_w570_v = ~(v_w2928_v & v_w2931_v);
	assign v_w6621_v = ~(v_w6592_v & v_w1003_v);
	assign v_w3709_v = ~(v_w3553_v & v_w3549_v);
	assign v_w3270_v = ~(v_w3126_v & v_w3269_v);
	assign v_w4689_v = ~(v_w4526_v | v_w4685_v);
	assign v_w2195_v = v_w48_v ^ v_w2163_v;
	assign v_w3111_v = ~(v_w2357_v & v_s429_v);
	assign v_w1258_v = ~(v_w1256_v & v_w1257_v);
	assign v_w6482_v = ~(v_w6472_v & v_w6471_v);
	assign v_w6820_v = ~(v_w6818_v | v_w6819_v);
	assign v_w976_v = ~(v_w1038_v & v_w1039_v);
	assign v_w5130_v = ~(v_w2416_v | v_w2370_v);
	assign v_w4960_v = ~(v_w2347_v & v_w2815_v);
	assign v_w2958_v = ~(v_s161_v & v_w564_v);
	assign v_w4281_v = v_w4277_v ^ v_w4280_v;
	assign v_w3527_v = ~(v_w2863_v & v_w2856_v);
	assign v_w1987_v = ~(v_w680_v & v_w1777_v);
	assign v_w465_v = ~(v_w6706_v & v_w6707_v);
	assign v_w1635_v = ~(v_w1052_v & v_s197_v);
	assign v_w5165_v = v_w5141_v & v_s27_v;
	assign v_w7568_v = ~(v_w608_v | v_w7081_v);
	assign v_w7096_v = ~(v_w7094_v | v_w7095_v);
	assign v_w8016_v = ~(v_s458_v ^ v_s378_v);
	assign v_w975_v = ~(v_in24_v ^ v_w1252_v);
	assign v_w4803_v = ~(v_w2448_v & v_w2791_v);
	assign v_w3267_v = ~(v_w3265_v & v_w3266_v);
	assign v_w3920_v = ~(v_w3912_v);
	assign v_w487_v = ~(v_w7655_v & v_w7656_v);
	assign v_w1107_v = ~(v_w1214_v & v_w850_v);
	assign v_w3310_v = ~(v_w3121_v | v_w2308_v);
	assign v_w2860_v = ~(v_w2839_v ^ v_w2859_v);
	assign v_w502_v = ~(v_w6610_v & v_w6615_v);
	assign v_w2894_v = ~(v_w2866_v | v_w2893_v);
	assign v_w1628_v = ~(v_w1249_v ^ v_w551_v);
	assign v_w4547_v = ~(v_w3527_v & v_w4546_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s446_v<=0;
	end
	else
	begin
	v_s446_v<=v_w499_v;
	end
	end
	assign v_w1414_v = ~(v_w1411_v | v_w1413_v);
	assign v_w6584_v = ~(v_s16_v & v_w562_v);
	assign v_w5624_v = ~(v_s267_v & v_w695_v);
	assign v_w3470_v = ~(v_w3452_v | v_w3469_v);
	assign v_w3635_v = ~(v_w3634_v & v_w3490_v);
	assign v_w1585_v = ~(v_w603_v | v_w1584_v);
	assign v_w8246_v = ~(v_w3517_v & v_w3519_v);
	assign v_w1546_v = ~(v_w1544_v & v_w1545_v);
	assign v_w5201_v = ~(v_w4326_v | v_w1_v);
	assign v_w294_v = ~(v_w5250_v & v_w5251_v);
	assign v_w7198_v = ~(v_s203_v & v_w7112_v);
	assign v_w5676_v = ~(v_s24_v & v_w695_v);
	assign v_w1431_v = ~(v_w666_v & v_s113_v);
	assign v_w1126_v = ~(v_w1125_v);
	assign v_w5546_v = ~(v_w5544_v & v_w5545_v);
	assign v_w2966_v = ~(v_w558_v & v_w2965_v);
	assign v_w156_v = v_s147_v & v_w5134_v;
	assign v_w5999_v = ~(v_s342_v & v_w528_v);
	assign v_w1038_v = ~(v_in26_v & v_w1258_v);
	assign v_w7683_v = ~(v_w7681_v | v_w7682_v);
	assign v_w2677_v = ~(v_w2478_v & v_w871_v);
	assign v_w4152_v = ~(v_w3412_v | v_w4151_v);
	assign v_w7857_v = ~(v_w651_v & v_w7678_v);
	assign v_w5338_v = ~(v_s228_v & v_w5293_v);
	assign v_w3726_v = ~(v_w3689_v & v_w3725_v);
	assign v_w6976_v = ~(v_w6972_v | v_w6975_v);
	assign v_w5241_v = ~(v_w2554_v | v_w1_v);
	assign v_w5646_v = ~(v_s120_v & v_w695_v);
	assign v_w2483_v = ~(v_w558_v & v_w2317_v);
	assign v_w3178_v = ~(v_w3177_v & v_w2639_v);
	assign v_w2289_v = v_s290_v ^ v_w2288_v;
	assign v_w6567_v = ~(v_w1052_v & v_s3_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s498_v<=0;
	end
	else
	begin
	v_s498_v<=v_w323_v;
	end
	end
	assign v_w5323_v = ~(v_w2601_v & v_w2309_v);
	assign v_w793_v = ~(v_w791_v | v_w792_v);
	assign v_w1838_v = ~(v_w607_v & v_w1837_v);
	assign v_w2479_v = ~(v_w2478_v & v_w2317_v);
	assign v_w7605_v = ~(v_w7603_v & v_w7604_v);
	assign v_w4786_v = ~(v_w674_v & v_s391_v);
	assign v_w2189_v = ~(v_w2177_v & v_w2188_v);
	assign v_w4149_v = v_w4145_v ^ v_w4148_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s385_v<=0;
	end
	else
	begin
	v_s385_v<=v_w433_v;
	end
	end
	assign v_w7576_v = ~(v_w1873_v | v_w7575_v);
	assign v_w5481_v = ~(v_w4863_v | v_w4692_v);
	assign v_w6763_v = ~(v_w1798_v & v_w1725_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s375_v<=0;
	end
	else
	begin
	v_s375_v<=v_w419_v;
	end
	end
	assign v_w6600_v = ~(v_w6599_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s62_v<=0;
	end
	else
	begin
	v_s62_v<=v_w70_v;
	end
	end
	assign v_w2053_v = ~(v_w1642_v & v_w2052_v);
	assign v_w4340_v = ~(v_w4338_v & v_w4339_v);
	assign v_w7827_v = ~(v_w654_v & v_w7826_v);
	assign v_w7225_v = ~(v_w7223_v | v_w7224_v);
	assign v_w7450_v = ~(v_w680_v | v_w919_v);
	assign v_w5604_v = ~(v_s41_v & v_w676_v);
	assign v_w4610_v = ~(v_w878_v & v_w4609_v);
	assign v_w7308_v = ~(v_w7306_v | v_w7307_v);
	assign v_w44_v = ~(v_w7899_v & v_w7900_v);
	assign v_w6502_v = ~(v_w664_v & v_s471_v);
	assign v_w2465_v = ~(v_w2463_v | v_w2464_v);
	assign v_w343_v = ~(v_w5638_v & v_w5639_v);
	assign v_w2050_v = ~(v_w2047_v & v_w1824_v);
	assign v_w7945_v = ~(v_s115_v & v_w2143_v);
	assign v_w651_v = v_w649_v & v_w650_v;
	assign v_w3574_v = ~(v_w1124_v);
	assign v_w6592_v = ~(v_w6579_v);
	assign v_w2654_v = v_w2653_v & v_s382_v;
	assign v_w3244_v = v_w2860_v | v_w2865_v;
	assign v_w367_v = ~(v_s504_v);
	assign v_w1212_v = ~(v_w612_v & v_s84_v);
	assign v_w6519_v = ~(v_w1701_v | v_w6518_v);
	assign v_w686_v = v_s85_v ^ v_w1780_v;
	assign v_w2764_v = ~(v_w2762_v & v_w2763_v);
	assign v_w6051_v = ~(v_w6050_v ^ v_s359_v);
	assign v_w5220_v = ~(v_w1646_v | v_w5145_v);
	assign v_w1001_v = ~(v_s29_v & v_w562_v);
	assign v_w2823_v = ~(v_w2822_v);
	assign v_w3321_v = ~(v_w2847_v | v_w2620_v);
	assign v_w5821_v = ~(v_w5819_v | v_w5820_v);
	assign v_w8208_v = ~(v_w5555_v & v_w5522_v);
	assign v_w5530_v = ~(v_w4524_v | v_w5123_v);
	assign v_w7144_v = v_s43_v & v_w7113_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s331_v<=0;
	end
	else
	begin
	v_s331_v<=v_w359_v;
	end
	end
	assign v_w7603_v = ~(v_w7602_v & v_w1685_v);
	assign v_w4538_v = ~(v_w3648_v & v_w4537_v);
	assign v_w6892_v = ~(v_w1096_v | v_w6579_v);
	assign v_w3480_v = ~(v_w3478_v & v_w3479_v);
	assign v_w4425_v = ~(v_w2343_v & v_w4424_v);
	assign v_w4275_v = ~(v_w3352_v & v_w4274_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s379_v<=0;
	end
	else
	begin
	v_s379_v<=v_w423_v;
	end
	end
	assign v_w7493_v = ~(v_w7325_v & v_w7492_v);
	assign v_w3023_v = ~(v_w3022_v ^ v_w3004_v);
	assign v_w2877_v = ~(v_s326_v | v_w2850_v);
	assign v_w186_v = ~(v_w5262_v & v_w5263_v);
	assign v_w4504_v = ~(v_w4451_v & v_w4503_v);
	assign v_w6151_v = ~(v_w5840_v & v_w6150_v);
	assign v_w563_v = v_w568_v & v_w612_v;
	assign v_w3860_v = ~(v_w3856_v & v_w3859_v);
	assign v_w4581_v = ~(v_w4580_v & v_w3604_v);
	assign v_w3559_v = ~(v_w3558_v);
	assign v_w1978_v = v_w1925_v & v_w1928_v;
	assign v_o4_v = v_w8045_v ^ v_w8055_v;
	assign v_w2048_v = v_w1824_v ^ v_w2047_v;
	assign v_w5111_v = ~(v_w5109_v & v_w5110_v);
	assign v_w3893_v = ~(v_w3891_v & v_w3892_v);
	assign v_w3898_v = ~(v_w3814_v & v_w3811_v);
	assign v_w1774_v = v_s96_v ^ v_w1773_v;
	assign v_w6710_v = ~(v_w6708_v & v_w6709_v);
	assign v_w3067_v = ~(v_w620_v | v_w3066_v);
	assign v_w5590_v = ~(v_s106_v & v_w676_v);
	assign v_w4880_v = v_s362_v & v_w674_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s387_v<=0;
	end
	else
	begin
	v_s387_v<=v_w435_v;
	end
	end
	assign v_w2494_v = ~(v_w2335_v | v_w617_v);
	assign v_w5023_v = ~(v_w5021_v | v_w5022_v);
	assign v_w6420_v = ~(v_w664_v & v_s468_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s438_v<=0;
	end
	else
	begin
	v_s438_v<=v_w490_v;
	end
	end
	assign v_w2542_v = ~(v_w2484_v & v_w2379_v);
	assign v_w2342_v = ~(v_w8214_v);
	assign v_w675_v = v_w5555_v;
	assign v_w8103_v = v_w1998_v | v_w2090_v;
	assign v_w1545_v = ~(v_w1051_v & v_s244_v);
	assign v_w7859_v = ~(v_w651_v & v_w7684_v);
	assign v_w3119_v = ~(v_w3109_v & v_w3118_v);
	assign v_w5044_v = ~(v_w5042_v & v_w5043_v);
	assign v_w3140_v = ~(v_s384_v & v_w1_v);
	assign v_w2113_v = ~(v_w2108_v | v_w2112_v);
	assign v_w5070_v = ~(v_w5068_v | v_w5069_v);
	assign v_w3679_v = ~(v_w3612_v | v_w3601_v);
	assign v_w7756_v = ~(v_w6842_v | v_w1919_v);
	assign v_w7134_v = ~(v_w7132_v | v_w7133_v);
	assign v_w1598_v = ~(v_w1500_v & v_w1597_v);
	assign v_w550_v = ~(v_w974_v | v_w975_v);
	assign v_w6887_v = ~(v_w6885_v | v_w6886_v);
	assign v_w2464_v = ~(v_w2429_v | v_w2417_v);
	assign v_w2660_v = v_s387_v ^ v_w2659_v;
	assign v_w7979_v = ~(v_s472_v & v_s392_v);
	assign v_w527_v = ~(v_w2143_v);
	assign v_w5093_v = ~(v_w2342_v | v_w5092_v);
	assign v_w1953_v = ~(v_w1951_v & v_w1952_v);
	assign v_w5043_v = ~(v_w2447_v & v_w2399_v);
	assign v_w5831_v = ~(v_w5829_v & v_w5830_v);
	assign v_w5944_v = ~(v_w892_v & v_w1342_v);
	assign v_w6480_v = ~(v_w6468_v | v_w6479_v);
	assign v_w4351_v = ~(v_w4054_v & v_s390_v);
	assign v_w1042_v = ~(v_in9_v ^ v_w1204_v);
	assign v_w5222_v = ~(v_w5220_v | v_w5221_v);
	assign v_w5807_v = ~(v_w5805_v | v_w5806_v);
	assign v_w7425_v = ~(v_w7418_v & v_w7424_v);
	assign v_w6350_v = ~(v_w1465_v | v_w6349_v);
	assign v_w7523_v = ~(v_w679_v | v_w1902_v);
	assign v_w2354_v = ~(v_w2352_v | v_w2353_v);
	assign v_w541_v = ~(v_w742_v & v_w743_v);
	assign v_w3988_v = ~(v_w756_v & v_w3735_v);
	assign v_w1694_v = ~(v_w1692_v & v_w1693_v);
	assign v_w4125_v = ~(v_w4115_v | v_w4124_v);
	assign v_w3946_v = ~(v_w3035_v | v_w3945_v);
	assign v_w2413_v = ~(v_s260_v & v_w697_v);
	assign v_w1967_v = ~(v_w1931_v | v_w1928_v);
	assign v_w2158_v = ~(v_s168_v | v_w2157_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s204_v<=0;
	end
	else
	begin
	v_s204_v<=v_w217_v;
	end
	end
	assign v_w7786_v = ~(v_w1919_v | v_w6744_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s508_v<=0;
	end
	else
	begin
	v_s508_v<=v_w386_v;
	end
	end
	assign v_w499_v = ~(v_w7834_v & v_w7835_v);
	assign v_w4335_v = ~(v_w4334_v & v_w690_v);
	assign v_w4719_v = ~(v_w4444_v & v_w3060_v);
	assign v_w524_v = ~(v_w6486_v & v_w6507_v);
	assign v_w5665_v = ~(v_w4082_v & v_w3060_v);
	assign v_w7717_v = ~(v_w654_v & v_w7716_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s146_v<=0;
	end
	else
	begin
	v_s146_v<=v_w155_v;
	end
	end
	assign v_w608_v = ~(v_w606_v | v_w607_v);
	assign v_w6348_v = ~(v_w657_v & v_s344_v);
	assign v_w7431_v = ~(v_w7394_v & v_w7430_v);
	assign v_w2521_v = ~(v_w2518_v & v_w2515_v);
	assign v_w383_v = ~(v_w5206_v & v_w5207_v);
	assign v_w1958_v = ~(v_s72_v | v_s71_v);
	assign v_w3584_v = ~(v_w3581_v & v_w3583_v);
	assign v_w495_v = ~(v_w7905_v & v_w7906_v);
	assign v_w4742_v = ~(v_w4526_v | v_w4741_v);
	assign v_w4406_v = ~(v_w825_v & v_w4405_v);
	assign v_w319_v = ~(v_w4152_v & v_w4168_v);
	assign v_w4078_v = ~(v_w690_v & v_w4077_v);
	assign v_w4570_v = ~(v_w3568_v & v_w4569_v);
	assign v_w5772_v = ~(v_s307_v & v_w529_v);
	assign v_w2982_v = ~(v_s115_v & v_w564_v);
	assign v_w7844_v = ~(v_w1783_v & v_w6585_v);
	assign v_w7541_v = ~(v_w7537_v | v_w7540_v);
	assign v_w2983_v = ~(v_w2779_v | v_w531_v);
	assign v_w3227_v = ~(v_s382_v & v_w1_v);
	assign v_w4493_v = ~(v_w2791_v | v_w968_v);
	assign v_w779_v = v_w1176_v & v_w1177_v;
	assign v_w25_v = ~(v_w5612_v & v_w5613_v);
	assign v_w6116_v = ~(v_w6114_v & v_w6115_v);
	assign v_w7069_v = ~(v_w7068_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s251_v<=0;
	end
	else
	begin
	v_s251_v<=v_w265_v;
	end
	end
	assign v_w5102_v = ~(v_w2369_v & v_w1131_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s86_v<=0;
	end
	else
	begin
	v_s86_v<=v_w94_v;
	end
	end
	assign v_w1347_v = ~(v_w1345_v & v_w1346_v);
	assign v_w6110_v = ~(v_w6108_v | v_w6109_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s358_v<=0;
	end
	else
	begin
	v_s358_v<=v_w397_v;
	end
	end
	assign v_w5980_v = ~(v_w662_v & v_w1026_v);
	assign v_w4932_v = ~(v_w674_v | v_w4931_v);
	assign v_w3226_v = ~(v_w2607_v & v_w2738_v);
	assign v_w7711_v = ~(v_w654_v & v_w7710_v);
	assign v_w6622_v = ~(v_w6620_v & v_w6621_v);
	assign v_w6689_v = ~(v_w6680_v & v_w6688_v);
	assign v_w8051_v = ~(v_w7979_v & v_w8050_v);
	assign v_w3712_v = ~(v_w3552_v & v_w3559_v);
	assign v_w519_v = ~(v_w6346_v & v_w6369_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s272_v<=0;
	end
	else
	begin
	v_s272_v<=v_w290_v;
	end
	end
	assign v_w3721_v = ~(v_w3596_v | v_w3720_v);
	assign v_w6357_v = ~(v_w6029_v | v_w6356_v);
	assign v_w2997_v = ~(v_w2995_v | v_w2996_v);
	assign v_w2392_v = ~(v_w2309_v | v_w2391_v);
	assign v_w4485_v = ~(v_w4483_v | v_w4484_v);
	assign v_w1034_v = ~(v_w1033_v | v_w899_v);
	assign v_w2211_v = ~(v_s128_v | v_s127_v);
	assign v_w6990_v = ~(v_s306_v & v_w656_v);
	assign v_w5096_v = ~(v_s260_v & v_w2347_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s369_v<=0;
	end
	else
	begin
	v_s369_v<=v_w412_v;
	end
	end
	assign v_w2725_v = v_w553_v ^ v_w2724_v;
	assign v_w6028_v = ~(v_w6026_v & v_w6027_v);
	assign v_w7765_v = ~(v_w7763_v & v_w7764_v);
	assign v_w1170_v = ~(v_w1169_v | v_s440_v);
	assign v_w4563_v = ~(v_w3559_v & v_w4562_v);
	assign v_w6742_v = ~(v_w6728_v | v_w6741_v);
	assign v_w5853_v = ~(v_w2137_v & v_w895_v);
	assign v_w336_v = ~(v_w3212_v & v_w3213_v);
	assign v_w4156_v = ~(v_w4145_v & v_w4148_v);
	assign v_w2265_v = ~(v_w2264_v);
	assign v_w1346_v = ~(v_w1052_v & v_s413_v);
	assign v_w7778_v = ~(v_w654_v & v_w7777_v);
	assign v_w4170_v = ~(v_w4169_v & v_w887_v);
	assign v_w373_v = ~(v_s505_v);
	assign v_w226_v = ~(v_w5636_v & v_w5637_v);
	assign v_w933_v = ~(v_w931_v | v_w932_v);
	assign v_w2218_v = ~(v_w2216_v & v_w2217_v);
	assign v_w5272_v = ~(v_w2343_v & v_w5271_v);
	assign v_w7900_v = ~(v_w651_v & v_w7807_v);
	assign v_w1960_v = ~(v_s46_v | v_w1959_v);
	assign v_w4397_v = ~(v_s425_v & v_w674_v);
	assign v_w4338_v = ~(v_w2985_v & v_w4319_v);
	assign v_w6910_v = ~(v_w6909_v | v_w953_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s377_v<=0;
	end
	else
	begin
	v_s377_v<=v_w421_v;
	end
	end
	assign v_w7536_v = ~(v_w680_v & v_w893_v);
	assign v_w7290_v = ~(v_w680_v | v_w1342_v);
	assign v_w2655_v = v_w2654_v & v_s383_v;
	assign v_w3478_v = ~(v_w3477_v & v_w2300_v);
	assign v_w1981_v = ~(v_w1976_v & v_w1980_v);
	assign v_w1137_v = ~(v_w2600_v);
	assign v_w720_v = v_w718_v & v_w719_v;
	assign v_w7889_v = ~(v_s102_v & v_w7876_v);
	assign v_w684_v = ~(v_w717_v & v_w28_v);
	assign v_w1786_v = ~(v_w657_v & v_w1190_v);
	assign v_w34_v = ~(v_s482_v);
	assign v_w1702_v = ~(v_w1374_v | v_w1701_v);
	assign v_w4424_v = v_w3468_v ^ v_w4423_v;
	assign v_w1936_v = ~(v_s66_v | v_s65_v);
	assign v_w1253_v = ~(v_s216_v & v_w1103_v);
	assign v_w5583_v = ~(v_w675_v & v_w5401_v);
	assign v_w2410_v = ~(v_w2357_v & v_s262_v);
	assign v_w1513_v = ~(v_w827_v | v_w8_v);
	assign v_w4331_v = ~(v_w2985_v & v_w4314_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s132_v<=0;
	end
	else
	begin
	v_s132_v<=v_w141_v;
	end
	end
	assign v_w2327_v = ~(v_w2326_v);
	assign v_w5176_v = ~(v_w693_v | v_w879_v);
	assign v_w3577_v = ~(v_w2738_v | v_w761_v);
	assign v_w7649_v = ~(v_w6011_v | v_w685_v);
	assign v_w4114_v = ~(v_w4056_v & v_s378_v);
	assign v_w3385_v = ~(v_w640_v & v_w2944_v);
	assign v_w4736_v = ~(v_w674_v & v_s397_v);
	assign v_w6808_v = ~(v_w1880_v ^ v_w6802_v);
	assign v_w5930_v = ~(v_w2117_v & v_w1866_v);
	assign v_w7128_v = ~(v_w1288_v | v_w7117_v);
	assign v_w1205_v = ~(v_s38_v & v_w1103_v);
	assign v_w5541_v = ~(v_w683_v & v_w5540_v);
	assign v_w3094_v = ~(v_w3092_v & v_w3093_v);
	assign v_w549_v = ~(v_in24_v | v_w1252_v);
	assign v_w2924_v = ~(v_w2358_v & v_s350_v);
	assign v_w521_v = ~(v_w6402_v & v_w6425_v);
	assign v_w1286_v = ~(v_w1282_v | v_w1285_v);
	assign v_w4172_v = ~(v_s311_v & v_w4056_v);
	assign v_w5311_v = ~(v_w5309_v | v_w5310_v);
	assign v_w42_v = ~(v_s484_v);
	assign v_w5289_v = ~(v_w2252_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s505_v<=0;
	end
	else
	begin
	v_s505_v<=v_w372_v;
	end
	end
	assign v_w7578_v = ~(v_w7576_v & v_w7577_v);
	assign v_w3055_v = ~(v_w3053_v & v_w3054_v);
	assign v_w6344_v = v_s195_v ^ v_w1465_v;
	assign v_w7527_v = ~(v_w7525_v & v_w7526_v);
	assign v_w3788_v = ~(v_w2980_v | v_w881_v);
	assign v_w4158_v = v_w4154_v ^ v_w4157_v;
	assign v_w7335_v = ~(v_w901_v | v_w680_v);
	assign v_w4020_v = ~(v_w4018_v | v_w4019_v);
	assign v_w3873_v = ~(v_w3848_v & v_w3851_v);
	assign v_w1182_v = ~(v_w1052_v & v_s13_v);
	assign v_w5441_v = ~(v_w5439_v | v_w5440_v);
	assign v_w8001_v = ~(v_s459_v | v_s295_v);
	assign v_w1617_v = ~(v_s323_v ^ v_w1153_v);
	assign v_w6440_v = v_w6433_v ^ v_w6439_v;
	assign v_w8253_v = ~(v_w608_v & v_w575_v);
	assign v_w4517_v = ~(v_w4515_v | v_w4516_v);
	assign v_w11_v = ~(v_w1992_v & v_w1994_v);
	assign v_w1996_v = ~(v_w1774_v & v_w882_v);
	assign v_w2690_v = ~(v_w2688_v & v_w2689_v);
	assign v_w3239_v = ~(v_w2607_v & v_w2910_v);
	assign v_w2661_v = ~(v_w2660_v & v_w2634_v);
	assign v_w6183_v = ~(v_w6181_v & v_w6182_v);
	assign v_w1852_v = ~(v_w1827_v | v_w1851_v);
	assign v_w6355_v = ~(v_w6353_v | v_w6354_v);
	assign v_w4703_v = ~(v_w2369_v & v_w3077_v);
	assign v_w3291_v = ~(v_w1016_v & v_w2639_v);
	assign v_w7708_v = ~(v_w765_v | v_w1782_v);
	assign v_w1569_v = ~(v_w1567_v | v_w1568_v);
	assign v_w5751_v = ~(v_w5749_v & v_w5750_v);
	assign v_w7209_v = ~(v_w7207_v | v_w7208_v);
	assign v_w2090_v = ~(v_w2088_v | v_w2089_v);
	assign v_w2662_v = ~(v_s387_v & v_w693_v);
	assign v_w7032_v = ~(v_w7030_v & v_w7031_v);
	assign v_w1697_v = ~(v_w870_v & v_w1696_v);
	assign v_w2772_v = ~(v_w2770_v & v_w2771_v);
	assign v_w2992_v = ~(v_w558_v & v_w2991_v);
	assign v_w3481_v = ~(v_w3476_v | v_w3480_v);
	assign v_w5083_v = ~(v_w2447_v & v_w2429_v);
	assign v_w2756_v = v_s111_v ^ v_w844_v;
	assign v_w3701_v = ~(v_w3529_v);
	assign v_w1540_v = v_w1374_v | v_w1539_v;
	assign v_w7721_v = ~(v_w7719_v | v_w7720_v);
	assign v_w4909_v = ~(v_w4908_v & v_w878_v);
	assign v_w7739_v = ~(v_w7737_v | v_w7738_v);
	assign v_w218_v = ~(v_w7872_v & v_w7873_v);
	assign v_w7122_v = ~(v_w7120_v | v_w7121_v);
	assign v_w4767_v = ~(v_w4766_v | v_w4589_v);
	assign v_w2577_v = ~(v_w2355_v & v_s221_v);
	assign v_w6867_v = ~(v_w656_v | v_w6866_v);
	assign v_w4955_v = ~(v_w4945_v & v_w4954_v);
	assign v_w7758_v = ~(v_w1783_v & v_w1437_v);
	assign v_w820_v = ~(v_w818_v & v_w819_v);
	assign v_w122_v = ~(v_w7760_v & v_w7761_v);
	assign v_w6964_v = ~(v_w6963_v & v_w6626_v);
	assign v_w3588_v = ~(v_w3142_v | v_w851_v);
	assign v_w5938_v = ~(v_w5936_v & v_w5937_v);
	assign v_w2671_v = ~(v_w2669_v & v_w2670_v);
	assign v_w4140_v = v_w4137_v ^ v_w4139_v;
	assign v_w3814_v = v_w3812_v | v_w3813_v;
	assign v_w1020_v = ~(v_w1070_v | v_w1071_v);
	assign v_w7553_v = v_w680_v | v_w7240_v;
	assign v_w3761_v = ~(v_w3735_v & v_w3060_v);
	assign v_w7623_v = ~(v_w1310_v | v_w7622_v);
	assign v_w6377_v = ~(v_w657_v & v_s345_v);
	assign v_w3187_v = ~(v_w2478_v & v_w963_v);
	assign v_w932_v = ~(v_w1373_v | v_w1883_v);
	assign v_w2239_v = ~(v_w8121_v);
	assign v_w6757_v = ~(v_s405_v & v_w656_v);
	assign v_w5911_v = ~(v_w662_v & v_w1813_v);
	assign v_w3463_v = ~(v_w3461_v & v_w3462_v);
	assign v_w4979_v = ~(v_w4977_v & v_w4978_v);
	assign v_w667_v = ~(v_w678_v ^ v_w19_v);
	assign v_w2562_v = ~(v_w2558_v);
	assign v_w3845_v = v_w3832_v | v_w3835_v;
	assign v_w5126_v = ~(v_w5125_v);
	assign v_w6619_v = ~(v_w934_v ^ v_w935_v);
	assign v_w1461_v = ~(v_w1458_v & v_w1460_v);
	assign v_w2754_v = ~(v_w2753_v | v_w557_v);
	assign v_w1419_v = ~(v_w1418_v | v_w1021_v);
	assign v_w1199_v = ~(v_s27_v & v_w1192_v);
	assign v_w4975_v = ~(v_w2369_v & v_w2833_v);
	assign v_w6473_v = ~(v_w6471_v ^ v_w6472_v);
	assign v_w3598_v = ~(v_w3596_v | v_w3597_v);
	assign v_w7674_v = ~(v_s358_v & v_w7667_v);
	assign v_w3719_v = ~(v_w3604_v & v_w3718_v);
	assign v_w7099_v = ~(v_w2126_v & v_w1837_v);
	assign v_w4671_v = ~(v_w4528_v | v_w4660_v);
	assign v_w5275_v = ~(v_w5273_v | v_w5274_v);
	assign v_w3494_v = ~(v_w2392_v);
	assign v_w7460_v = ~(v_w679_v | v_w1823_v);
	assign v_w4699_v = ~(v_w8218_v);
	assign v_w6276_v = ~(v_w6241_v & v_w6244_v);
	assign v_w1110_v = v_w8102_v ^ v_keyinput_27_v;
	assign v_w2280_v = ~(v_s111_v | v_w2168_v);
	assign v_w7783_v = ~(v_w6773_v & v_w7782_v);
	assign v_w2039_v = ~(v_w2033_v);
	assign v_w4729_v = ~(v_w4727_v & v_w4728_v);
	assign v_w5577_v = ~(v_w675_v & v_w5376_v);
	assign v_w4902_v = ~(v_w4900_v & v_w4901_v);
	assign v_w3457_v = ~(v_s8_v & v_w1192_v);
	assign v_w876_v = ~(v_w2241_v & v_w880_v);
	assign v_w2640_v = ~(v_w2639_v & v_w2575_v);
	assign v_w641_v = ~(v_w2013_v | v_w2029_v);
	assign v_w2543_v = ~(v_w558_v & v_w2297_v);
	assign v_w5041_v = v_w2442_v ^ v_w2438_v;
	assign v_w1498_v = ~(v_w1495_v | v_w1497_v);
	assign v_w3941_v = ~(v_w3563_v);
	assign v_w7608_v = ~(v_w1419_v | v_w7607_v);
	assign v_w6031_v = ~(v_w42_v | v_w889_v);
	assign v_w6083_v = ~(v_w6076_v & v_w6082_v);
	assign v_w7616_v = ~(v_w1352_v & v_w1364_v);
	assign v_w6371_v = ~(v_w6361_v & v_w6360_v);
	assign v_w7589_v = ~(v_w7253_v ^ v_w6585_v);
	assign v_w7750_v = ~(v_w1919_v | v_w6859_v);
	assign v_w1410_v = ~(v_w875_v & v_s406_v);
	assign v_w6712_v = ~(v_w6711_v & v_w6626_v);
	assign v_w2349_v = ~(v_w2344_v & v_w2348_v);
	assign v_w7292_v = ~(v_w7290_v | v_w7291_v);
	assign v_w3407_v = ~(v_w3403_v | v_w3406_v);
	assign v_w6470_v = ~(v_s114_v & v_w6429_v);
	assign v_w3578_v = ~(v_w3577_v);
	assign v_w1494_v = ~(v_w874_v & v_s306_v);
	assign v_w3644_v = v_w8114_v ^ v_keyinput_37_v;
	assign v_w4550_v = ~(v_w4535_v | v_w4549_v);
	assign v_w5615_v = ~(v_w675_v & v_w5540_v);
	assign v_w7388_v = ~(v_w680_v | v_w831_v);
	assign v_w4874_v = ~(v_w4872_v | v_w4873_v);
	assign v_w5475_v = ~(v_w5473_v | v_w5474_v);
	assign v_w4871_v = ~(v_w2369_v & v_w2993_v);
	assign v_w7695_v = ~(v_w834_v | v_w1782_v);
	assign v_w2954_v = ~(v_s364_v & v_w2358_v);
	assign v_w2921_v = ~(v_w2919_v & v_w2920_v);
	assign v_w5630_v = ~(v_s232_v & v_w695_v);
	assign v_w4079_v = ~(v_w4054_v & v_s377_v);
	assign v_w1637_v = ~(v_w1635_v & v_w1636_v);
	assign v_w7846_v = ~(v_w654_v & v_w7845_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s168_v<=0;
	end
	else
	begin
	v_s168_v<=v_w178_v;
	end
	end
	assign v_w7594_v = ~(v_w1769_v & v_w1761_v);
	assign v_w4184_v = ~(v_w4182_v & v_w4183_v);
	assign v_w2182_v = ~(v_s169_v | v_w2171_v);
	assign v_w7584_v = ~(v_w6659_v | v_w7583_v);
	assign v_w6252_v = ~(v_s215_v & v_w888_v);
	assign v_w666_v = v_w665_v;
	assign v_w1829_v = ~(v_w1828_v & v_w989_v);
	assign v_w1799_v = ~(v_s12_v & v_w1374_v);
	assign v_w532_v = ~(v_w7235_v & v_w7236_v);
	assign v_w6489_v = ~(v_w6487_v & v_w6488_v);
	assign v_w991_v = ~(v_w990_v | v_w531_v);
	assign v_w1443_v = v_w969_v ^ v_w796_v;
	assign v_w6337_v = ~(v_w6018_v | v_w1644_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s40_v<=0;
	end
	else
	begin
	v_s40_v<=v_w47_v;
	end
	end
	assign v_w7443_v = ~(v_w687_v | v_w839_v);
	assign v_w4027_v = ~(v_w4026_v & v_w2233_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s306_v<=0;
	end
	else
	begin
	v_s306_v<=v_w329_v;
	end
	end
	assign v_w1005_v = ~(v_s34_v & v_w562_v);
	assign v_w459_v = ~(v_w4679_v & v_w4694_v);
	assign v_w4415_v = ~(v_w851_v | v_w4414_v);
	assign v_w2491_v = ~(v_w2489_v | v_w2490_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s471_v<=0;
	end
	else
	begin
	v_s471_v<=v_w524_v;
	end
	end
	assign v_w7867_v = ~(v_w651_v & v_w7710_v);
	assign v_w5216_v = ~(v_w693_v | v_w2929_v);
	assign v_w986_v = ~(v_w984_v | v_w985_v);
	assign v_w8240_v = ~(v_w6908_v | v_w6920_v);
	assign v_w3957_v = ~(v_w3950_v | v_w3956_v);
	assign v_w5810_v = ~(v_w826_v | v_w633_v);
	assign v_w3952_v = ~(v_w3035_v | v_w3731_v);
	assign v_w3058_v = ~(v_w3055_v | v_w3057_v);
	assign v_w7848_v = ~(v_w1783_v & v_w7636_v);
	assign v_w3639_v = ~(v_w3536_v | v_w3531_v);
	assign v_w5483_v = ~(v_w5481_v | v_w5482_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s517_v<=0;
	end
	else
	begin
	v_s517_v<=v_w483_v;
	end
	end
	assign v_w4488_v = ~(v_w4486_v | v_w4487_v);
	assign v_w7112_v = ~(v_w612_v | v_s475_v);
	assign v_w5240_v = ~(v_w1506_v | v_w5145_v);
	assign v_w7469_v = ~(v_w7462_v & v_w7459_v);
	assign v_w3680_v = ~(v_w3678_v & v_w3679_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s314_v<=0;
	end
	else
	begin
	v_s314_v<=v_w339_v;
	end
	end
	assign v_w4474_v = ~(v_w3647_v | v_w4473_v);
	assign v_w6424_v = v_w8109_v ^ v_keyinput_33_v;
	assign v_w4115_v = ~(v_w3312_v & v_w4114_v);
	assign v_w718_v = ~(v_w721_v | v_s320_v);
	assign v_w5400_v = ~(v_w5398_v | v_w5399_v);
	assign v_w4994_v = ~(v_w2261_v | v_w2581_v);
	assign v_w3914_v = ~(v_w3913_v & v_w1017_v);
	assign v_w7675_v = ~(v_w7068_v | v_w1919_v);
	assign v_w5014_v = ~(v_w2363_v | v_w2261_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s244_v<=0;
	end
	else
	begin
	v_s244_v<=v_w257_v;
	end
	end
	assign v_w2752_v = ~(v_w2750_v & v_w2751_v);
	assign v_w1147_v = ~(v_w1145_v | v_w1146_v);
	assign v_w750_v = ~(v_w591_v | v_w752_v);
	assign v_w7899_v = ~(v_s37_v & v_w7876_v);
	assign v_w5733_v = ~(v_w892_v & v_w917_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s476_v<=0;
	end
	else
	begin
	v_s476_v<=v_w530_v;
	end
	end
	assign v_w6885_v = ~(v_w656_v | v_w6884_v);
	assign v_w3280_v = ~(v_w2391_v | v_w2606_v);
	assign v_w5603_v = ~(v_w5555_v & v_w5486_v);
	assign v_w468_v = ~(v_w7821_v & v_w7822_v);
	assign v_w2801_v = ~(v_w2795_v | v_w2800_v);
	assign v_w456_v = ~(v_w4699_v & v_w4714_v);
	assign v_w2988_v = ~(v_w2981_v | v_w2987_v);
	assign v_w4181_v = v_s299_v ^ v_w4169_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s24_v<=0;
	end
	else
	begin
	v_s24_v<=v_w26_v;
	end
	end
	assign v_w7535_v = ~(v_w687_v & v_w1187_v);
	assign v_w4831_v = ~(v_w4829_v | v_w4830_v);
	assign v_w2766_v = v_w404_v ^ v_w2648_v;
	assign v_w7949_v = ~(v_s110_v & v_w2143_v);
	assign v_w6574_v = ~(v_w1976_v & v_w1991_v);
	assign v_w4884_v = ~(v_w4882_v & v_w4883_v);
	assign v_w5914_v = ~(v_w5912_v | v_w5913_v);
	assign v_w4315_v = ~(v_w2984_v ^ v_w4314_v);
	assign v_w2876_v = ~(v_s123_v & v_w565_v);
	assign v_w6217_v = ~(v_w6215_v & v_w6216_v);
	assign v_w5894_v = ~(v_w5890_v | v_w5893_v);
	assign v_w4057_v = ~(v_s263_v & v_w4056_v);
	assign v_w6230_v = ~(v_w6029_v | v_w6229_v);
	assign v_w6284_v = ~(v_w6282_v | v_w6283_v);
	assign v_w5677_v = ~(v_w4082_v & v_w3118_v);
	assign v_w8173_v = v_w3373_v & v_w1139_v;
	assign v_w8045_v = ~(v_w7985_v | v_w8044_v);
	assign v_w6874_v = v_w1865_v ^ v_w6870_v;
	assign v_w6749_v = ~(v_w6745_v & v_w758_v);
	assign v_w5785_v = ~(v_w5783_v & v_w5784_v);
	assign v_w7362_v = ~(v_w1642_v | v_w680_v);
	assign v_w3110_v = ~(v_w593_v & v_s23_v);
	assign v_w4730_v = ~(v_w4526_v | v_w4725_v);
	assign v_w5663_v = ~(v_w4082_v & v_w2722_v);
	assign v_w5767_v = ~(v_w1073_v ^ v_w5766_v);
	assign v_w1612_v = ~(v_w1606_v | v_w839_v);
	assign v_w2201_v = ~(v_s147_v | v_s146_v);
	assign v_w1728_v = ~(v_w797_v);
	assign v_w2191_v = ~(v_w2189_v & v_w2190_v);
	assign v_w1754_v = ~(v_w666_v & v_s418_v);
	assign v_w2331_v = v_w2328_v & v_w1034_v;
	assign v_w894_v = ~(v_w1999_v ^ v_w1075_v);
	assign v_w5277_v = ~(v_w2458_v & v_w5276_v);
	assign v_w3492_v = ~(v_w825_v | v_w2890_v);
	assign v_w656_v = ~(v_w655_v);
	assign v_w4276_v = ~(v_s363_v & v_w4056_v);
	assign v_w4579_v = ~(v_w4577_v | v_w4578_v);
	assign v_w2070_v = ~(v_w2068_v & v_w2069_v);
	assign v_w702_v = ~(v_in32_v & v_w545_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s32_v<=0;
	end
	else
	begin
	v_s32_v<=v_w36_v;
	end
	end
	assign v_w5726_v = ~(v_w662_v & v_w1350_v);
	assign v_w3810_v = ~(v_w2856_v | v_w3735_v);
	assign v_w358_v = ~(v_w4234_v & v_w4240_v);
	assign v_w404_v = ~(v_s511_v);
	assign v_w4319_v = ~(v_w8126_v);
	assign v_w6154_v = ~(v_w6152_v & v_w6153_v);
	assign v_w3647_v = ~(v_w3528_v | v_w3532_v);
	assign v_w4740_v = ~(v_w4738_v | v_w4739_v);
	assign v_w1792_v = ~(v_w875_v & v_s452_v);
	assign v_w939_v = v_w2676_v & v_w2680_v;
	assign v_w7718_v = ~(v_s214_v & v_w7667_v);
	assign v_w4271_v = ~(v_w4264_v & v_w4270_v);
	assign v_w4988_v = ~(v_w4987_v & v_w673_v);
	assign v_w2872_v = ~(v_w2358_v & v_s362_v);
	assign v_w7053_v = ~(v_w7051_v & v_w7052_v);
	assign v_w586_v = v_w2893_v | v_w2948_v;
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s207_v<=0;
	end
	else
	begin
	v_s207_v<=v_w220_v;
	end
	end
	assign v_w6878_v = ~(v_w1798_v & v_w1453_v);
	assign v_w2237_v = ~(v_w2236_v | v_w531_v);
	assign v_w4787_v = ~(v_w3005_v & v_w2347_v);
	assign v_w5209_v = ~(v_w1443_v | v_w5145_v);
	assign v_w3118_v = ~(v_w3116_v & v_w3117_v);
	assign v_w4364_v = ~(v_w4348_v | v_w4346_v);
	assign v_w7961_v = ~(v_s38_v & v_w2143_v);
	assign v_w508_v = ~(v_w6059_v & v_w6067_v);
	assign v_w6250_v = ~(v_w6228_v & v_w6226_v);
	assign v_w1793_v = ~(v_w1791_v & v_w1792_v);
	assign v_w6397_v = ~(v_s345_v & v_w6373_v);
	assign v_w6315_v = ~(v_w6305_v & v_w6304_v);
	assign v_w7622_v = ~(v_w1312_v | v_w7621_v);
	assign v_w1369_v = ~(v_w1366_v & v_w1368_v);
	assign v_w4848_v = v_w4488_v ^ v_w4457_v;
	assign v_w3212_v = ~(v_w3210_v | v_w3211_v);
	assign v_w6114_v = ~(v_s244_v & v_w889_v);
	assign v_w4235_v = ~(v_w2851_v ^ v_s202_v);
	assign v_w1174_v = ~(v_w943_v | v_w1173_v);
	assign v_w1664_v = ~(v_w1239_v ^ v_w751_v);
	assign v_w4001_v = ~(v_w3995_v & v_w4000_v);
	assign v_w578_v = ~(v_w576_v & v_w577_v);
	assign v_w5291_v = ~(v_s167_v & v_w5134_v);
	assign v_w1662_v = ~(v_w1659_v & v_w1661_v);
	assign v_w2590_v = ~(v_w2575_v);
	assign v_w2346_v = v_s292_v ^ v_w2345_v;
	assign v_w7954_v = ~(v_w527_v & v_w1813_v);
	assign v_w3306_v = ~(v_w3304_v & v_w3305_v);
	assign v_w6049_v = ~(v_w1579_v | v_w6048_v);
	assign v_w4088_v = ~(v_w4086_v | v_w4087_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s97_v<=0;
	end
	else
	begin
	v_s97_v<=v_w105_v;
	end
	end
	assign v_w1048_v = ~(v_w1046_v & v_w1047_v);
	assign v_w1992_v = ~(v_w1923_v & v_w651_v);
	assign v_w2883_v = ~(v_s124_v ^ v_w2882_v);
	assign v_w7165_v = ~(v_w7163_v | v_w7164_v);
	assign v_w5408_v = ~(v_w5405_v & v_w5407_v);
	assign v_w888_v = ~(v_w657_v);
	assign v_w5729_v = ~(v_w5727_v | v_w5728_v);
	assign v_w401_v = ~(v_s510_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s309_v<=0;
	end
	else
	begin
	v_s309_v<=v_w332_v;
	end
	end
	assign v_w5178_v = ~(v_w5176_v | v_w5177_v);
	assign v_w1812_v = ~(v_w1363_v & v_w1729_v);
	assign v_w1003_v = ~(v_w1001_v & v_w1002_v);
	assign v_w5290_v = ~(v_w2248_v | v_s174_v);
	assign v_w5039_v = ~(v_w880_v | v_w5038_v);
	assign v_w3354_v = ~(v_w3352_v & v_w3353_v);
	assign v_w5943_v = ~(v_w5941_v | v_w5942_v);
	assign v_w5018_v = ~(v_w5017_v | v_w4526_v);
	assign v_w6155_v = v_w1514_v ^ v_w6154_v;
	assign v_w1072_v = v_w599_v | v_w2065_v;
	assign v_w2172_v = ~(v_s166_v | v_w2171_v);
	assign v_w8061_v = ~(v_w7995_v | v_w7996_v);
	assign v_w38_v = ~(v_w5672_v & v_w5673_v);
	assign v_w7153_v = ~(v_w7151_v | v_w7152_v);
	assign v_w4636_v = ~(v_w4444_v & v_w2671_v);
	assign v_w5085_v = ~(v_w2465_v ^ v_w2460_v);
	assign v_w2637_v = ~(v_w2623_v | v_w2636_v);
	assign v_w86_v = ~(v_w5664_v & v_w5665_v);
	assign v_w4280_v = ~(v_w4278_v & v_w4279_v);
	assign v_w5526_v = ~(v_w964_v | v_w2602_v);
	assign v_w6043_v = ~(v_w6020_v & v_w6042_v);
	assign v_w2925_v = ~(v_w2923_v & v_w2924_v);
	assign v_w5690_v = ~(v_w892_v & v_w766_v);
	assign v_w4567_v = ~(v_w4566_v | v_w3633_v);
	assign v_w6538_v = ~(v_w6537_v & v_w6516_v);
	assign v_w5482_v = ~(v_w3574_v | v_w2602_v);
	assign v_w2949_v = ~(v_w699_v & v_s176_v);
	assign v_w7457_v = ~(v_w687_v & v_w1823_v);
	assign v_w6696_v = ~(v_w1788_v & v_w1350_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s393_v<=0;
	end
	else
	begin
	v_s393_v<=v_w442_v;
	end
	end
	assign v_w3769_v = ~(v_w760_v & v_w881_v);
	assign v_w4314_v = ~(v_w4312_v | v_w4313_v);
	assign v_w3728_v = ~(v_w3470_v | v_w3727_v);
	assign v_w4195_v = ~(v_w3205_v | v_w4194_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s479_v<=0;
	end
	else
	begin
	v_s479_v<=v_w7_v;
	end
	end
	assign v_w3008_v = ~(v_w3006_v & v_w3007_v);
	assign v_w6581_v = ~(v_w6577_v | v_w6580_v);
	assign v_w4546_v = ~(v_w3647_v & v_w4545_v);
	assign v_w5399_v = ~(v_w4863_v | v_w4885_v);
	assign v_w7477_v = ~(v_w7341_v & v_w7476_v);
	assign v_w3591_v = ~(v_w3576_v | v_w3590_v);
	assign v_w2019_v = ~(v_w723_v ^ v_w536_v);
	assign v_w7656_v = ~(v_w1975_v & v_w1972_v);
	assign v_w8226_v = ~(v_w1298_v & v_w1750_v);
	assign v_w1983_v = ~(v_w1963_v | v_w1982_v);
	assign v_w1736_v = ~(v_w1352_v & v_w1735_v);
	assign v_w3742_v = ~(v_w3737_v & v_w3740_v);
	assign v_w3004_v = ~(v_w2765_v | v_w3003_v);
	assign v_w8136_v = v_w2319_v | v_w2323_v;
	assign v_w408_v = ~(v_w4308_v & v_w4309_v);
	assign v_w2139_v = ~(v_w1761_v | v_w2138_v);
	assign v_w1183_v = ~(v_w874_v & v_s449_v);
	assign v_w2000_v = ~(v_w1999_v ^ v_w1067_v);
	assign v_w908_v = v_w906_v & v_w907_v;
	assign v_w6917_v = ~(v_w6915_v ^ v_w6916_v);
	assign v_w751_v = ~(v_w749_v | v_w750_v);
	assign v_w52_v = ~(v_w7145_v & v_w7146_v);
	assign v_w5699_v = ~(v_w662_v & v_w1297_v);
	assign v_w3670_v = ~(v_w3633_v | v_w3669_v);
	assign v_w1471_v = ~(v_w1126_v | v_w1096_v);
	assign v_w5215_v = ~(v_s123_v & v_w5141_v);
	assign v_w6394_v = ~(v_w6389_v & v_w6393_v);
	assign v_w6836_v = ~(v_w6834_v | v_w6835_v);
	assign v_w4138_v = ~(v_s239_v & v_w4116_v);
	assign v_w5877_v = ~(v_w2137_v & v_w1026_v);
	assign v_w5586_v = ~(v_s117_v & v_w676_v);
	assign v_w3822_v = v_w3818_v | v_w3821_v;
	assign v_w6903_v = ~(v_w6901_v | v_w6902_v);
	assign v_w5817_v = ~(v_s438_v & v_w529_v);
	assign v_w4588_v = ~(v_w2457_v | v_w880_v);
	assign v_w64_v = v_s56_v & v_w7107_v;
	assign v_w5910_v = ~(v_s404_v & v_w528_v);
	assign v_w4274_v = ~(v_w2884_v & v_w887_v);
	assign v_w6677_v = ~(v_w6675_v | v_w6676_v);
	assign v_w2011_v = ~(v_w723_v ^ v_w989_v);
	assign v_w315_v = ~(v_w2637_v & v_w2640_v);
	assign v_w1075_v = ~(v_w1074_v);
	assign v_w5650_v = ~(v_s112_v & v_w695_v);
	assign v_w2145_v = ~(v_w181_v & v_w2144_v);
	assign v_w4205_v = ~(v_w4054_v & v_s317_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s252_v<=0;
	end
	else
	begin
	v_s252_v<=v_w267_v;
	end
	end
	assign v_w1101_v = ~(v_w1100_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s461_v<=0;
	end
	else
	begin
	v_s461_v<=v_w514_v;
	end
	end
	assign v_w8066_v = v_w8065_v ^ v_keyinput_2_v;
	assign v_w8129_v = ~(v_w6527_v & v_w6528_v);
	assign v_w7706_v = v_w6978_v ^ v_keyinput_30_v;
	assign v_w169_v = ~(v_w7881_v & v_w7882_v);
	assign v_w1575_v = v_w608_v | v_w575_v;
	assign v_w6830_v = ~(v_w6641_v & v_w6829_v);
	assign v_w7310_v = ~(v_w7305_v & v_w7308_v);
	assign v_w3384_v = v_w639_v & v_w3244_v;
	assign v_w2018_v = v_w2017_v & v_w729_v;
	assign v_w1095_v = ~(v_w1469_v & v_w1470_v);
	assign v_w3133_v = ~(v_w3127_v & v_w3132_v);
	assign v_w3805_v = ~(v_w2926_v | v_w881_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s478_v<=0;
	end
	else
	begin
	v_s478_v<=v_w1_v;
	end
	end
	assign v_w78_v = v_s70_v & v_w7107_v;
	assign v_w6811_v = ~(v_w6809_v & v_w6810_v);
	assign v_w6980_v = ~(v_w1787_v & v_w788_v);
	assign v_w6722_v = ~(v_w656_v | v_w6721_v);
	assign v_w4507_v = ~(v_w4505_v | v_w4506_v);
	assign v_w7152_v = v_w7112_v & v_s84_v;
	assign v_w2181_v = ~(v_s166_v | v_w2174_v);
	assign v_w452_v = ~(v_w4721_v & v_w4735_v);
	assign v_w1912_v = ~(v_w1911_v ^ v_w859_v);
	assign v_w1660_v = ~(v_w1125_v | v_w1095_v);
	assign v_w5682_v = ~(v_s6_v & v_w695_v);
	assign v_w6816_v = ~(v_w656_v | v_w6815_v);
	assign v_w7777_v = ~(v_w7775_v & v_w7776_v);
	assign v_w1337_v = ~(v_w1335_v & v_w1336_v);
	assign v_w6495_v = ~(v_w6029_v | v_w6494_v);
	assign v_w4377_v = ~(v_w690_v & v_w4376_v);
	assign v_w6324_v = ~(v_w657_v & v_s338_v);
	assign v_w5725_v = ~(v_s411_v & v_w528_v);
	assign v_w196_v = ~(v_w5462_v & v_w5471_v);
	assign v_w5077_v = ~(v_w2347_v & v_s261_v);
	assign v_w1331_v = ~(v_w1330_v | v_w1180_v);
	assign v_w7273_v = ~(v_w687_v & v_w1067_v);
	assign v_w2867_v = ~(v_w699_v & v_s175_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s388_v<=0;
	end
	else
	begin
	v_s388_v<=v_w436_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s417_v<=0;
	end
	else
	begin
	v_s417_v<=v_w468_v;
	end
	end
	assign v_w1325_v = ~(v_w1066_v & v_w1324_v);
	assign v_w4991_v = ~(v_w4989_v & v_w4990_v);
	assign v_w7561_v = ~(v_w647_v | v_w1028_v);
	assign v_w569_v = ~(v_w568_v);
	assign v_w7086_v = ~(v_w7084_v & v_w7085_v);
	assign v_w5940_v = ~(v_w5938_v | v_w5939_v);
	assign v_w7028_v = ~(v_w7024_v & v_w7027_v);
	assign v_w6531_v = ~(v_w6021_v | v_w6530_v);
	assign v_w1502_v = v_w587_v & v_s7_v;
	assign v_w5515_v = ~(v_w683_v & v_w5514_v);
	assign v_w941_v = ~(v_w8107_v);
	assign v_w1057_v = ~(v_w1055_v | v_w1056_v);
	assign v_w4345_v = ~(v_w4336_v | v_w4344_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s105_v<=0;
	end
	else
	begin
	v_s105_v<=v_w113_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s436_v<=0;
	end
	else
	begin
	v_s436_v<=v_w488_v;
	end
	end
	assign v_w4443_v = ~(v_w4441_v | v_w4442_v);
	assign v_w6055_v = v_w8073_v ^ v_keyinput_9_v;
	assign v_w372_v = ~(v_w5716_v & v_w5722_v);
	assign v_w3727_v = ~(v_w3687_v & v_w3726_v);
	assign v_w1824_v = ~(v_w1624_v);
	assign v_w1354_v = v_w850_v ^ v_w1214_v;
	assign v_w6267_v = ~(v_w6251_v | v_w6255_v);
	assign v_w4270_v = ~(v_w4269_v & v_w692_v);
	assign v_w7127_v = ~(v_w7118_v & v_w1277_v);
	assign v_w6071_v = ~(v_w6053_v);
	assign v_w6795_v = ~(v_w6791_v & v_w6794_v);
	assign v_w349_v = ~(v_w5737_v & v_w5745_v);
	assign v_w4489_v = ~(v_w4457_v | v_w4488_v);
	assign v_w4664_v = ~(v_w4663_v & v_w673_v);
	assign v_w4532_v = ~(v_w4531_v & v_w2341_v);
	assign v_w7689_v = v_w7687_v & v_w7688_v;
	assign v_w6932_v = v_w1858_v ^ v_w6912_v;
	assign v_w8029_v = ~(v_w8027_v | v_w8028_v);
	assign v_w7137_v = v_w7113_v & v_s431_v;
	assign v_w2672_v = ~(v_w872_v | v_w2606_v);
	assign v_w694_v = ~(v_w604_v & v_w2194_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s395_v<=0;
	end
	else
	begin
	v_s395_v<=v_w444_v;
	end
	end
	assign v_w7911_v = ~(v_s9_v & v_w7876_v);
	assign v_w5974_v = ~(v_w5970_v | v_w5973_v);
	assign v_w8084_v = ~(v_w937_v ^ v_w552_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s13_v<=0;
	end
	else
	begin
	v_s13_v<=v_w14_v;
	end
	end
	assign v_w136_v = v_s127_v & v_w5134_v;
	assign v_w1336_v = ~(v_w666_v & v_s415_v);
	assign v_w318_v = ~(v_w5015_v & v_w5033_v);
	assign v_w1247_v = ~(v_w612_v & v_s203_v);
	assign v_w1679_v = ~(v_w1094_v & v_w1678_v);
	assign v_w4011_v = ~(v_w3687_v & v_w4010_v);
	assign v_w7876_v = ~(v_w651_v);
	assign v_w3562_v = ~(v_w864_v | v_w3025_v);
	assign v_w6761_v = ~(v_w6759_v | v_w6760_v);
	assign v_w7147_v = ~(v_w1781_v | v_w529_v);
	assign v_o14_v = ~(v_w8021_v ^ v_w8022_v);
	assign v_w4242_v = ~(v_w4235_v & v_w4238_v);
	assign v_w8056_v = ~(v_w7985_v | v_w7986_v);
	assign v_w6935_v = ~(v_w6911_v ^ v_w6912_v);
	assign v_w1810_v = ~(v_w1323_v | v_w1066_v);
	assign v_w3402_v = ~(v_w3401_v & v_w1139_v);
	assign v_w1450_v = ~(v_w1448_v & v_w1449_v);
	assign v_w2138_v = ~(v_w2137_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s6_v<=0;
	end
	else
	begin
	v_s6_v<=v_w6_v;
	end
	end
	assign v_w7145_v = ~(v_w6012_v | v_w7144_v);
	assign v_w5652_v = ~(v_s373_v & v_w695_v);
	assign v_w5826_v = ~(v_w1302_v | v_w2135_v);
	assign v_w5567_v = ~(v_w675_v & v_w5336_v);
	assign v_w2121_v = ~(v_w1970_v & v_w1990_v);
	assign v_w4135_v = ~(v_w4056_v & v_s295_v);
	assign v_w6341_v = ~(v_w1644_v & v_w6316_v);
	assign v_w2023_v = v_w602_v ^ v_w2017_v;
	assign v_w2670_v = ~(v_w2355_v & v_s33_v);
	assign v_w6320_v = ~(v_w1626_v & v_w6298_v);
	assign v_w7898_v = ~(v_w651_v & v_w7801_v);
	assign v_w3642_v = v_w8070_v ^ v_keyinput_5_v;
	assign v_w6229_v = ~(v_w6226_v ^ v_w6228_v);
	assign v_w715_v = ~(v_w714_v | v_s302_v);
	assign v_w7331_v = ~(v_w1436_v | v_w680_v);
	assign v_w4891_v = ~(v_w4890_v & v_w878_v);
	assign v_w4701_v = ~(v_w4700_v & v_w878_v);
	assign v_w1509_v = ~(v_w1051_v & v_s226_v);
	assign v_w1940_v = ~(v_w1934_v & v_w1939_v);
	assign v_w3961_v = ~(v_w3342_v | v_w3731_v);
	assign v_w5426_v = ~(v_s179_v & v_w5386_v);
	assign v_w956_v = ~(v_w2967_v & v_w1088_v);
	assign v_w2217_v = ~(v_s142_v | v_s140_v);
	assign v_w4408_v = ~(v_w1083_v & v_w4407_v);
	assign v_w2537_v = ~(v_w2378_v | v_w557_v);
	assign v_w5392_v = ~(v_w5390_v | v_w5391_v);
	assign v_w880_v = ~(v_w866_v);
	assign v_w1941_v = ~(v_s58_v | v_s57_v);
	assign v_w2424_v = ~(v_w698_v & v_s257_v);
	assign v_w341_v = ~(v_w4964_v & v_w4974_v);
	assign v_w8206_v = v_w4619_v & v_w4620_v;
	assign v_w7253_v = ~(v_w1796_v);
	assign v_w7078_v = ~(v_w7074_v | v_w7077_v);
	assign v_w6978_v = v_w1596_v ^ v_w980_v;
	assign v_w6467_v = ~(v_w6464_v ^ v_w6466_v);
	assign v_w538_v = ~(v_w537_v);
	assign v_w1727_v = ~(v_w1714_v | v_w799_v);
	assign v_w108_v = ~(v_w7161_v & v_w7162_v);
	assign v_w6806_v = ~(v_w6592_v & v_w1817_v);
	assign v_w4934_v = ~(v_w2342_v | v_w4933_v);
	assign v_w2269_v = ~(v_s218_v | v_w2268_v);
	assign v_w4746_v = ~(v_w2448_v & v_w3338_v);
	assign v_w6104_v = ~(v_w6102_v & v_w6103_v);
	assign v_w3359_v = ~(v_w2893_v | v_w2941_v);
	assign v_w7291_v = ~(v_w687_v | v_w1350_v);
	assign v_w4598_v = ~(v_w4596_v | v_w4597_v);
	assign v_w3886_v = ~(v_w3882_v & v_w3885_v);
	assign v_w6568_v = ~(v_w1758_v & v_w6567_v);
	assign v_w5195_v = ~(v_s103_v & v_w5141_v);
	assign v_w2084_v = ~(v_w1337_v | v_w2083_v);
	assign v_w6098_v = ~(v_w6096_v & v_w6097_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s428_v<=0;
	end
	else
	begin
	v_s428_v<=v_w479_v;
	end
	end
	assign v_w5504_v = ~(v_w4642_v | v_w5123_v);
	assign v_w7447_v = ~(v_w687_v | v_w920_v);
	assign v_w3522_v = ~(v_w3521_v | v_w2618_v);
	assign v_w7548_v = ~(v_w7252_v | v_w7256_v);
	assign v_w7178_v = ~(v_s112_v & v_w7113_v);
	assign v_w7546_v = ~(v_w7544_v | v_w7545_v);
	assign v_w6943_v = ~(v_s324_v & v_w656_v);
	assign v_w6164_v = ~(v_w6157_v & v_w6163_v);
	assign v_w2047_v = v_w1999_v ^ v_w1632_v;
	assign v_w1006_v = ~(v_w756_v | v_w2690_v);
	assign v_w2822_v = v_s312_v ^ v_w2796_v;
	assign v_w5027_v = ~(v_w5016_v & v_w5026_v);
	assign v_w4544_v = ~(v_w3646_v | v_w4543_v);
	assign v_w5103_v = ~(v_w5101_v & v_w5102_v);
	assign v_w2358_v = v_w2357_v;
	assign v_w1666_v = ~(v_w1665_v | v_w8_v);
	assign v_w6132_v = ~(v_w1539_v & v_w6104_v);
	assign v_w3779_v = ~(v_w881_v | v_w968_v);
	assign v_w1580_v = ~(v_w1579_v);
	assign v_w7806_v = ~(v_w1783_v & v_w917_v);
	assign v_w6297_v = ~(v_w657_v & v_s324_v);
	assign v_w7615_v = ~(v_w1731_v | v_w7614_v);
	assign v_w2468_v = ~(v_w2466_v | v_w2467_v);
	assign v_w4911_v = ~(v_w4909_v & v_w4910_v);
	assign v_w8237_v = ~(v_w3369_v | v_w2620_v);
	assign v_w7635_v = ~(v_w7594_v & v_w7634_v);
	assign v_w7237_v = ~(v_w6569_v);
	assign v_w3344_v = ~(v_w3341_v | v_w3343_v);
	assign v_w3081_v = ~(v_w3068_v | v_w3080_v);
	assign v_w1236_v = ~(v_s123_v & v_w1192_v);
	assign v_w1691_v = ~(v_w1402_v | v_w1690_v);
	assign v_w5322_v = ~(v_s238_v & v_w5293_v);
	assign v_w7057_v = ~(v_w2127_v | v_w566_v);
	assign v_w6204_v = ~(v_w6029_v | v_w6203_v);
	assign v_w2306_v = ~(v_w2304_v | v_w2305_v);
	assign v_w727_v = ~(v_w2011_v | v_w788_v);
	assign v_w2510_v = ~(v_w2504_v | v_w2500_v);
	assign v_w1078_v = v_w8097_v ^ v_keyinput_24_v;
	assign v_w6308_v = ~(v_w664_v & v_s464_v);
	assign v_w2683_v = ~(v_w2355_v & v_s39_v);
	assign v_w277_v = ~(v_w3399_v & v_w3400_v);
	assign v_w5378_v = ~(v_s199_v & v_w5293_v);
	assign v_w4311_v = ~(v_w3441_v & v_w4310_v);
	assign v_w665_v = ~(v_w668_v | v_w669_v);
	assign v_w1084_v = ~(v_w2785_v & v_w2786_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s115_v<=0;
	end
	else
	begin
	v_s115_v<=v_w124_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s5_v<=0;
	end
	else
	begin
	v_s5_v<=v_w5_v;
	end
	end
	assign v_w3128_v = ~(v_s1_v | v_w401_v);
	assign v_w1856_v = ~(v_w1606_v);
	assign v_w6376_v = ~(v_s122_v & v_w888_v);
	assign v_w7268_v = ~(v_w7266_v & v_w7267_v);
	assign v_w8134_v = v_w1287_v ^ v_w2097_v;
	assign v_w4505_v = ~(v_w782_v | v_w4504_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s63_v<=0;
	end
	else
	begin
	v_s63_v<=v_w71_v;
	end
	end
	assign v_w1343_v = v_w461_v ^ v_w1165_v;
	assign v_w7125_v = v_w7112_v & v_s24_v;
	assign v_w5128_v = ~(v_w2428_v | v_w3495_v);
	assign v_w2761_v = ~(v_w2753_v);
	assign v_w2248_v = ~(v_w2247_v);
	assign v_w7755_v = ~(v_s159_v & v_w7742_v);
	assign v_w1374_v = v_w672_v;
	assign v_w872_v = ~(v_w2671_v);
	assign v_w529_v = ~(v_s519_v);
	assign v_w307_v = ~(v_w5846_v & v_w5851_v);
	assign v_w1466_v = ~(v_w1374_v | v_w1465_v);
	assign v_w4606_v = ~(v_w4603_v | v_w4605_v);
	assign v_w3357_v = ~(v_w3244_v & v_w638_v);
	assign v_w6019_v = ~(v_w6018_v);
	assign v_w2817_v = ~(v_s209_v & v_w699_v);
	assign v_w8044_v = ~(v_w7986_v | v_w8043_v);
	assign v_w1599_v = ~(v_w1052_v & v_s207_v);
	assign v_w4087_v = ~(v_w3336_v | v_w691_v);
	assign v_w245_v = ~(v_w5630_v & v_w5631_v);
	assign v_w2357_v = v_w592_v & v_w544_v;
	assign v_w5433_v = ~(v_w683_v & v_w5432_v);
	assign v_w6459_v = ~(v_w6456_v ^ v_w6458_v);
	assign v_w994_v = v_in17_v ^ v_w1229_v;
	assign v_w1902_v = ~(v_w1297_v);
	assign v_w921_v = ~(v_w1134_v | v_w920_v);
	assign v_w7164_v = ~(v_w7117_v | v_w1703_v);
	assign v_w3431_v = ~(v_w3430_v & v_w1139_v);
	assign v_w2776_v = ~(v_w2775_v & v_w2152_v);
	assign v_w613_v = ~(v_w671_v);
	assign v_w1281_v = ~(v_w870_v & v_w1280_v);
	assign v_w1000_v = ~(v_w757_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s444_v<=0;
	end
	else
	begin
	v_s444_v<=v_w496_v;
	end
	end
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s56_v<=0;
	end
	else
	begin
	v_s56_v<=v_w64_v;
	end
	end
	assign v_w4452_v = ~(v_w3561_v | v_w3566_v);
	assign v_w6741_v = ~(v_w656_v | v_w6740_v);
	assign v_w1440_v = v_s367_v ^ v_w1421_v;
	assign v_w491_v = ~(v_w6658_v & v_w6672_v);
	assign v_w2508_v = ~(v_w2506_v & v_w2507_v);
	assign v_w1145_v = ~(v_w6590_v & v_w6572_v);
	assign v_w1683_v = ~(v_w1682_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s405_v<=0;
	end
	else
	begin
	v_s405_v<=v_w454_v;
	end
	end
	assign v_w1307_v = ~(v_w1303_v | v_w1306_v);
	assign v_w2732_v = ~(v_w2358_v & v_s397_v);
	assign v_w4250_v = ~(v_w4249_v & v_w4231_v);
	assign v_w6680_v = ~(v_w6679_v & v_w884_v);
	assign v_w6636_v = ~(v_w6634_v & v_w6635_v);
	assign v_w4450_v = ~(v_w852_v & v_w3142_v);
	assign v_w1726_v = ~(v_w1725_v);
	assign v_w1254_v = ~(v_w612_v & v_s213_v);
	assign v_w3029_v = ~(v_w2358_v & v_s394_v);
	assign v_w347_v = ~(v_w5894_v & v_w5901_v);
	assign v_w1734_v = ~(v_w1342_v);
	assign v_w5498_v = ~(v_s186_v & v_w5293_v);
	assign v_w1387_v = ~(v_s107_v & v_w562_v);
	assign v_w929_v = ~(v_w1818_v | v_w1880_v);
	assign v_w5648_v = ~(v_s366_v & v_w695_v);
	assign v_w6608_v = ~(v_w1787_v);
	assign v_w1210_v = ~(v_w1208_v & v_w1209_v);
	assign v_w12_v = ~(v_w7973_v & v_w7974_v);
	assign v_w2204_v = ~(v_s151_v | v_s150_v);
	assign v_w3047_v = ~(v_w8066_v);
	assign v_w7193_v = ~(v_w7191_v | v_w7192_v);
	assign v_w1473_v = v_w714_v & v_s7_v;
	assign v_w8123_v = v_w8122_v ^ v_keyinput_42_v;
	assign v_w7098_v = ~(v_s158_v & v_w1140_v);
	assign v_w2294_v = v_w2293_v;
	assign v_w3879_v = v_w3839_v | v_w3842_v;
	assign v_w7771_v = ~(v_w6815_v & v_w7770_v);
	assign v_w935_v = ~(v_w8227_v);
	assign v_w8002_v = ~(v_s458_v | v_s378_v);
	assign v_w8097_v = ~(v_w1076_v | v_w1077_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s121_v<=0;
	end
	else
	begin
	v_s121_v<=v_w130_v;
	end
	end
	assign v_w5194_v = ~(v_w5192_v | v_w5193_v);
	assign v_w3449_v = v_w3447_v & v_w3448_v;
	assign v_w8243_v = v_w8242_v ^ v_keyinput_121_v;
	assign v_w4272_v = ~(v_w2929_v | v_w4041_v);
	assign v_w6442_v = ~(v_s341_v & v_w6399_v);
	assign v_w5092_v = v_w2326_v ^ v_w2336_v;
	assign v_w1105_v = ~(v_in14_v & v_w1220_v);
	assign v_w5032_v = ~(v_w2342_v | v_w5031_v);
	always@(posedge v_in1_v )
	begin
	if(reset)
	begin
	v_s102_v<=0;
	end
	else
	begin
	v_s102_v<=v_w110_v;
	end
	end
	assign v_w410_v = ~(v_w7181_v & v_w7182_v);
	assign v_w4666_v = ~(v_w2265_v & v_w753_v);
	assign v_w8161_v = v_w8160_v ^ v_keyinput_67_v;
	assign v_w6888_v = ~(v_s345_v & v_w656_v);
	assign v_w2945_v = ~(v_w2944_v);
	assign v_w6596_v = ~(v_w6595_v & v_w757_v);
	assign v_w1164_v = v_w1163_v | v_s404_v;
	assign v_w7136_v = ~(v_w528_v | v_w1931_v);
	assign v_w7686_v = ~(v_s243_v & v_w7667_v);
	assign v_w6940_v = ~(v_w1140_v & v_w1617_v);
	assign v_w4766_v = v_w4499_v ^ v_w4452_v;
	assign v_w4679_v = ~(v_w4677_v | v_w4678_v);
	assign v_w5239_v = ~(v_s309_v & v_w5140_v);
	assign v_w4625_v = v_w3630_v ^ v_w4517_v;
	assign v_w2449_v = ~(v_w2448_v & v_w2439_v);
	assign v_w1701_v = ~(v_w1700_v);
	assign v_w1018_v = ~(v_in18_v & v_w1232_v);
	assign v_w3378_v = ~(v_w3376_v | v_w3377_v);
	assign v_w522_v = ~(v_w6431_v & v_w6453_v);
	assign v_w4704_v = ~(v_w4702_v & v_w4703_v);
	assign v_w6454_v = ~(v_w1424_v & v_w6444_v);
	assign v_w258_v = ~(v_w7679_v & v_w7680_v);
	assign v_w7047_v = v_w1548_v ^ v_w1587_v;
	assign v_w4918_v = ~(v_w4916_v & v_w4917_v);
	assign v_w5140_v = ~(v_w1192_v | v_s1_v);
	assign v_w2893_v = ~(v_w2888_v | v_w2892_v);
	assign v_w4490_v = ~(v_w2993_v | v_w2991_v);
	assign v_w185_v = ~(v_s489_v);
	assign v_w6298_v = ~(v_w6296_v & v_w6297_v);
	assign v_w1570_v = ~(v_w665_v & v_s356_v);
	assign v_w2390_v = ~(v_w2388_v & v_w2389_v);
endmodule
